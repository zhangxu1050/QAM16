��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O �ٝ�l�������V��fE��v�-�Q��Rj&	ڭE�����<��1`5��o"�l�&��3J���m\�tu*&W�N[��H��j	�����[6ҊZq]ս"�!z���z��r5����nk�/�v����~��8r��,��:ƛ���M-$��e�~4=#�g�L�C�� \3˂��M�~���Wξ���G��Iǎ�S��IhU�_J]��;'M�J�ӕk�g��b��v��ҵ푣�~���/O�ׅ���08n2�B�
|Rh�ώX�T`;<�/y��m�=q;a�߸h�{���ð�t���f��
*tLb?�S
n�Uj�
�J ~���lAoT?�!d$��1�-;�59�C@YO*��x6S�����0��*�?��'d�>�fCŝ�ug��ENm�HKj���i�@�����&�F�kZ�8���E���b,>�#z��Ƭu?�_ͥ-�BH�k>�K
 ���AS���+�����>�E�c��?$�*rJ>&+a�#PS\�-����r�٭|�!��S����7�9���[|)���
�;>(i�>����Z;C��>��T���:1x��L;Utu�S׫E���.�ޒ12�Ꮠ���Z��|�*Wټ �iVr�+��<wzl����d:�:w�"����:Z
�Μ���IU���~�w�HJ��P����#�>����2��Ms��_�'����~J<!�
?V�9�o���bM��0��� �E��S��k�[�s�L�O��WX��-3B��O�
+ʮj��"O��P~���Q�_����~�����ؽ��̍ϲ�=��e��I�n1Rn�YDy|�/�\��v]A�>����M���z�v�s+�a/G��TB�w4xnРCҪd�����iV�sB�郡�1Z��������0~��,K��|(�{�| B��\
)����b`�j>j�O�
��6����|z5&~萤�h�����Gq�/�!�`�'仁"0�q3�X L ��+ ��_�-I�<��ܯ����F.G��C<NdĨoÝ��F*�T����PE��<r�5��^��E�Jd?@	I���/HRd�X� 7��z�t���M����d�
Ƴ�%���[v2�5%$\=� 2����G6ȥ�+� ����s��@*����"�%s�I ��CP�[@��3�\��:��  �1�p��\������yє��+O� ��a	��6�;��<Y;/(~gT�� �^�cL�~���f��N�dmy�C����$�ѱ �Qկ��1��Ͼ&aA�y�;&�Ӟkw�]⬆[$���qgG����}�>h��&zo��*�J[���T��Tq��U�SvB� C~1�e,��>�+��I��E^�0��B��Q(�;�Q���zR��|���eRD�iv*��z�T<���}hܶ��F��t93FgMl)�"�u�>�]�b����st���▸(��Q��L���wDY�4h��c�Ӛd�h����g�2vl��ҋ�m��f3��áV孳��(9�]C�N�*}� �a�e]���� q~�y۳��@2X9�#O�<A�S�٘���3�eyPB�2���>�v�J7SN2�2�Fǁ37pc�t{��|�����(�p�ymO1���h6���<k�;�{��h�p�sq�6�8zxдÄLi�;�K�[����ä́-��\�5k#|&5u�b1�R�xN*h$)y���[w�Uԍs�����b|m�C:%�'1T �6
��Oq�_�"6�1a=Н�\lf\QQ�)By{��֬gf[�Ͼ&N�����L���u�\�t�̦ѐ��5�!�TB���gcp��7�C����~��"�!ÍF����=�P\��.���4�:z���⯝��&^w�6˴����0۽�X������:�S��j��E��3Sz���Z-A�0�7)-�#��N�����*1/F(5�-��+�V�*T�c�ԭk�n���U �l�0��~�1��w[M��93e�Ͳ�o>EKQs��P���8����9װ^�>��f�Yy����;&Z�ݻ�=�� s�D����*
J@�3A{���
p:Thw��4,[&�,�O��+�p��d�z>{��ל(w`�S���{��WR��V-Sd�M��O�H"� }���U%��^���u�]k��#�Fd$�\&��*�Dc��B�%���}-2�EO�&��Z�N}sb�,��]R\��d�Iݞ=���H7�Gijc��}����sd'��x �Y�K�IZv�uU���k&�C#(�{�'�v�S�������@\�����oJ7����6m7�@m��s�F!@BD��p��)q* R0���m���j�{k_ ���EA��E�c��Hr��3'F��)�(o�c&��:���1K��8p��^K�9Bԯ���AsX�])A�k���r��l-��q��Rl���K�i��0+n���&}�{����f~q�}f��5�-�!ݭ�i9r?!(�R(�{����yr��k"b��>yQ�T�x��zz1�M-��N�usB�R��f9��>��Z�$���LRl�59v��B<e�$JQ^�dO1���_�����nt,H���z��P��d��"p��~��3Jis܋?N޼���ę�=ǎY��tm(�q�|ٷ�����g�\~��KA{Ѯ��ǆB;�<����0;��͈�I�y~���ڎ�3����������)�eR�sq�TB�aA��BQPkզuu���\r�[�bG�_�m�<$�Fz}��/�m�L���re�a��KM��y ��;���Y]@��o�s��\P]�W �1)���S/6��k$�c�Ɛ��n&��?�6�h�x>Ik����3-Kױ?V@�L���R.���=�[�ڊy«=���&��a����4�y��B��׎XƉ��S��\����V�gd�:B��콩ٲ�?d`�qf��Y��Rg�F&A��M�/���+a�>��k���{��>�D
y	O7��g�Χ�N�e{=�ku�um,.����E�'�i��}���]|,n�07������u��0��)��͵�9q/����SE>֦-�������EwYs�$:K�2E(������O��ЛD���$�=#^��hd���睅��6�f���Ƥ���Գ� qO��ec��������<���eYK�9#��$��\��
��v+?܊�B������AH-����W�/�12���:��"U�.þ3rx)C��1�!�w��!�Fm�ɐx�Q�d,�������NT�.���FC�tA�U���k��/�u��:$<~�P�n!r@8ܔ�i���Do����4<q������B$���qBZ�mB����{N-9�?m�����C�s.H����L�_�`��ː�yU�G�b�N���v��>��&��)a�ʅ���V� s4�1	Os0mV)�)xp�H�t�Ĵ��Hq[GV{ৱ�k<Wq�Yչ��Q#�YZ?����^��g�}��(WyN%�J+����$4~S��R�h����-v�J0�$�*bv�!�eZ��� ����t4�"���3��22K���~����:��/r�a֨$���\R�;����ܜU{�w�w)Ы����5���t ���)z��Y8����iA޲ YBATW߮=��k�2��i-����k?��������� KX����f�
�9�}8\*?�] �yɸ�>��4��?3�e�MpN�{��e�����u��+ӑ���b�̰� 
i� &����\I��;�=5
E#K(2�ME2�o�X������^d4�/݉b��H"c���]껼��]�8!�9����2��_�pyx�,J�Y� ��w������Z�k�w���R'�}�,�7�['���܋�dޘ�C]J����^R?�v�DZ�z�Bd�TQ�
=��g�ڲo���0��D~&�'A��
���ߧ2�i�����z�XA���/\��L�:EE�o˻MW>�������)��	�:�7�'C0!+~Ǧ�hu�$MJA]+4�ǳL[K��E�V�����K��7H)��O3��}jK��7���g�c���d#ՋcLj�*���5yN��{<-4K�m;U�\�&1N��-Q�_�����20�l��N:*cv���G8��	��{��r%�4e�ċZ-������$�����W!����D�zA#���5�]���R�B�^�w�[����m�"�b��T�Q�q�wC�,���e����|.��V�oXL�0O"�ea��+��H�O *������=뽲[�Lħw2�`�
�#^��
f�g�H2\�v�>��Lq.���q��Lr }
HCҟ���c�3=p�~F�nTb5?�������� ]����w�$,n�賬�Fe.��)��I6�����S �=����U����h��t��8Hh|=���l-7�/�0*�:�G���{�D��QL���;ֶ� |�ۋ��c�͌��1|��µd\�3 �,��H�pd��1m�ÆD��ws�qn�E�z>�Wf�4J�5�P���l� a��)�5���p�a��F��;ᘣ�Â��'M��a�0]�����p7��ϸ@h���i4�Ȧ)�����6[<�Ԡsȁ�3��e�p7h�&/W�^��*����Wl�����+�܏`�N##匃�k�.��f_�g�u��T�{h��ΠlV�3i�U�����"O5�׽��q$�a�(�8�>P��UT`vY��4�i��n��&j����:��9�|�"���e҂���n�8�(��l@9iF^���C)]���K+��?�`G�#;l�0�FxZ;V�٘?,�=�]�X�hG箶92A��,ֆ��������s.7����������M�J�0"��N|A3�*��pH�Q�b�?����b�#�2���j��͵������)C�㻵�{
lSվz���A�3sw�"k	)�J��������Eg�v�d�4Vd�s�f�(�����֫^1��؎.�����/^6$��>ۘ�d!�O���Ð���+`V������ᖒN8��VVz��u�t���?(���a�ߘש���#���bsx<+߶C���W������b6*d�>bS�8��S�R~E����&����l&�h����I� r(��$�p|�nU����7�!��diZ���=�M
D�K*P6{$��m�����U�v���b>"�Y�.u賧��H��<�R��S�K��g��Qb>��_t'����B�y[c��b���"f΢�=I��EÚ�2/gG�dv�)�vO�U8��x���YGէ��$TfI?���+3p�܏���n 2;�&d3���y(�vw,堭��8�����g�q���쟒@�9������#��/�t���h�4�����R~�t�HYۧ��[Pi�ǚ������!�!e��A�Pn-� (ߜ�k9s� �M�L(�a���M�A�1�1��C�ƚ�ArLo�{�c���{l��א�kco�8_�H��s�����g)����*J� �`I:?��gCuhbd��j�W���A9;L�H���x�y�����+�� ����!��#�ۙoI���-��_G��
pF�xS��<��߈>�s��W��HJ��{��-�b#���+6����jUI ��Ú�5�E�"�f�wȝ' ڿK�&u���x��HJ��@��� S�ܸ����k��2�Y3r�S��=|ċ����6j'+������i)P����+c���ӄ��X�j��*�Y\���E�|R�;�G��	5D���Ο�8���6���'��^:�~��Q�f�+�{L:�3�?�J�8
jO|yl�'C#}6�^�����]�Xq0��ae�D���ܐ��������b���I�_�BM�.4��s�1f8w3eҬ`�g�z��wjm�V�#c��g���~R=N�;��'{\��i������+�`T��#��fb��wtd2vSs��J�0�0A�uѐlO�n 0�4�]	�P2:+0o+Q\M�{sa@�<� ��ʵ,Yk�5�+�#�&�(�kـNe�	�m��yv7������j���k���ϸ��1�>-Ti���S'�� �S�73�M�ރ\�౿��s��1�;Mh�2j�~��v�(���������
�{�^�I��x��l�w�/�������Il;�\G�8z��Rߩ<p|U-���}�[v��:�DoC�#.�SNƯ"@N2�_��`���=�}��Z{���ⷤMb��(`����y֢j.��7��Bo��|NP�8Ew?��#��N���M�c/>|�
zo��W��龎C���ٰM�JĖTV����q�ּ�d9p��uGQ/:V��o�����s1;����rH�־6>:�`��;������Ƈ dY� ��w�X��_x(�[NǺ"��iګ�؎���KN6��z��Z���)�~Q�}.z�,�ƚ���q��c���XJ���9���� �ײWa�&�ϖGq�=HW��<��_�����Q�UʄW&r ���i�K�#�̈́�,��\��0=1��ܻ�����B�'�]Asno��.#BC�Ez�|�k�}Y���*��+�]W��zy�L����@�	Q�?��?�;6��綟��,�=u[�]��j����<ɞK��C���L�����2�Ti��]������<�K�@����e�U��;����vC0��v�zϕ�vO��pف�?��@gc�Ssm?�&u�(�H��?Riԏ���iE�ݠ�/���AE���w�q��7���"/W�_-�HR�u_��!P"k�+NI�������b��ű��_ZU�:FQ���u=<]��U��(�e�H����n[Z������oS�X�ǳ�o�#�|�5��8v|� ���X`y���w�$d8=1iZ��`L���i����'��?���9~ o�ǡ"�����х�E�!k6�Nc�G�")�W�8�!�*@�D�P����x~b-��B���OT��S���}���F��dÞ�~���֬7�}*�[���/�"In����4��Fj��������tf��?�y�A2�J>-������BVF��T�n��@���y�y=�Ю�/P