��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��W N��|C��#�N' ���x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`h��>��ׯ�=>)m��U���T���딣0&_���X0���2|	p��rw@	@us�犢����g��	K���yq�`݊�|���"rG�
���}�\���V�S/+��K��������طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-�!�5�?�����?9S��m�S� ���������	x]�m�Je{q�Я�mڍ'T����X澗�)�$���:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA�����h1�t��⫓���RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|?_W�\I��^�َ2V�N�u�k1i�f1?�نN��_�Q�L���E#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l������ ���yX�,I\�Z˻r���V�>!�/�7��u���nEA�i�+���6�Pr"?D2BC��5��Yk"1/���%	v3�.�z,yri�y�!�3]o��in�m��+Ȑ E�������?9���Z=%�l8������t�iZ]XF�������̘�иܖ��i (LW4WɆ&6�\]�4�6�t���]7K�6�á�~O�Y-�E�f��Z�>)��`�U+�PA����Kp&�@���k�փ��㛋��X���`��wl��h�ٙ���O����
��j��3�_� ��"����5'C��[���ԍ�7�"�����=���aˤ�� �e>����C8�����G%�MP3�u��N�v{�ҋX������S8�J�]=��R�^Ƒ����"X��[��Q[R�7�⒍~���u��N�v{�ҋX������S8�J�]=��R�^Ƒ����"X��[�d�a�4$�[�л���7��|g�Y�'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<��/�^�Ӭ����
L'���Xw s4S�'�i��иܖ��%����8��T�\ ��P�%.^F�	��lC��U�T�\ ��+�_0c �.�wK��� �ҋX����>��l%i�-�Aɀ��{l�f|�ό���.��_F�k-�7Ê7�E�4'���Xw����������)ҵ��]�!����M[��Ǣ����K? T�ҋX����*�QN��� ]���f�+��T��/o��إP�e`b�T=am���� F���9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8����W N��|C��ɹ���� �v���:�5����`K�aVD�C��l"�u<�rם4�S��ł�!r��Z����p�U���o氶�#7�V��hW
l�L��M�,���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9��
�����B�E`^n�&�
_�n�@/%{�;����Q��ǺΕ�f�f3'�g��U-�e���b P_�F�����CY���<�;�L���9��Xv7�j�i���TR�^Ƒ�ӽ�}^v��Z鎬�������(���`$�P.eE���lC��U�T�\ ��y�.�`L⯣�v[����_��ƕW��V�6IWJE�$��dg0J/��=��K�E��{#6�ae�ˑ���CY���<����,D/�Ú6��css2�����y:�u�J�@����gG��l��`�����C�#�,Z鎬�������(���P����ˮ��lC��U�T�\ ��i3�|)sՀ�6�S2v"Ohƪڈm�d�٣��c�A�L'R�o�����5�%]���a(􆿳���2����.��DP֞ -o�Ild�:�n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u��ArV�~ ��ç�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gG�[bGf���`M��
��
��D&e�2l��4�i�2�X&l����_::���`y����@����gG���:qJӰe4I��
��D&e�2l��4�i�2�X&l����H�^=�h{&|#9���b!��u�+�uB;y��TB	6е��*ܑe�W����n�4����ԻV8����ei��"X��[�d�a�4$�e�0
A���̹U�����r���	w	Qrk)�7JS�����,MLG򬉢��S��ȍry��	��yso6L�4��'��v��@�������>[HÛON�?��!�`�(i3,ԯ���gn��Ab�%^��}Dq�f��N�v�1�c����L�{�E����F�Z�>)�ώ�~+�ݗ�r'Z1p8��e�j�!�`�(i3,ԯ���gn�J����� ��}Dq�f��.��Ԕ�	���ZX�E����F���8�TP��IL;��$��8_�8���&�'�al��p�I�PD�na"�,�>E��4];ˍH����TI��Ԫ,щ�"��Wʁ�Wp7�:�!�`�(i3x�]�V���t�����[F�a�+�ީ�%��Wp7�:�!�`�(i37�ܥ��2�`e7��9��×�>���`�)J*~���f��0�5tU���D	��U�l>o��|���bǬ�=��I(�c��U��j�fH��>d]=]A��O�T=�4e=��-Y�VN�=��7p�J��PWV����ft���}�k�����5	��{�OF8F���m¡�����hWK{m35%7� ��yDgx�]�V���t���CՐ3��F<Y��j3��� Q�N��*���������@�%�I=�4e=��-V�׍A�ž_�F���yso6L%+�&��v��@�������>[HNl����!�`�(i3�E����F�Z�>)�ώ�~+�ݗ����>[H����&?�!�`�(i3�E����F�Z�>)�ώ�~+�ݗ�r'Z1p8��Y"H���!�`�(i3�E����F�Z�>)�����˟y� �>��|���;��x��B5��E����F���8�TPm=_g}b��t��6�5�p���PF��W�!�`�(i3зq8�Ј)w�<�_N��M��+?���C&����Wʁ�w�*�fBg�!�`�(i3���+�J��U<o^.K�}�{��$&XT
��"{phDJ��3Y� 2��4����7
!�`�(i37�ܥ��2�`e7��9��×�>��� �>��|~���f�A�������E����F���8�TP��@E�`�8���&�Q�$_��^�|n�M�!�`�(i3=]A��O�T=�4e=��-"w߻Y��}Dq�f���R�㺺|:=�C��Z��N�l������l>o��|���JLm|�Q'݀�=���SCh��{<qH�~�!�`�(i37�ܥ��2���kܪ���*�LNm�t����}ꇐ�622���k˗S�d�!�`�(i3x�]�V���t�����[F�a�+����ܗ�J���z!����k˗S�d�зq8�Ј)w�<�_N`E�cvR+��}Dq�f��v1a{J��]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=��I(�c��U��j��k˗S�d�"�,�>E��4];ˍH����TI��Ԫ,щ�"��<H��(����O��B�r�������5	��{�OF8F���m¡�����hWK{m35%,�!�H<Ȳ��+�J��U<o^.K�}qW8+����8���&�qr�^*4y-X��;^��J1!be�=]A��O�T=�4e=��-V�׍A���}Dq�f���*����	��Y��71{!�`�(i3���D	��U�l>o��|��b��7u�� л�b����\�TfZ!4Я\�rƛ�}�ٸW�{vK &�k+���!�`�(i3!�`�(i3=]A��O�T=�4e=��-�z�)lq���a���8���&�1籢��N�o!�`�(i3!�`�(i3�����5	��{�OF8�_�/�ߥ$Nx���t��y(�����������(������%�G"QL�)w�<�_N�eب�-�t���k��-��Wf<��;����7�/>�"�Ax!�`�(i3!�`�(i3x�]�V��;���Ӧ��Gjh�rO-�����`J�^���gJ!�`�(i3!�`�(i3�E����F���8�TPT֟��B�:УWKŃ����`J�*���u�Ww3i�|�!�`�(i3�E����F���8�TPT֟��B�:УWKŃz�q�����GO����!�`�(i3!�`�(i3�E����F�Z�>)�����˟y�u3v��U�DnK�]_!C6%K�pıN�c뵣�"�,�>E��4];ˍH�,t����t�&Fc$�n}��]"danS����˥����AB9���w�!�`�(i3x�]�V���T�3�R��	���I����r����$^�y1�\GD@�F��qW��Ґ�Yj���|��1��$�V��b�s������=���aI���;E�@%���8�a�"��FX1��t��L̿��$|�/|�z)�_m-�oq��f�}������!H�P|�����7JS�����,MLG�	�6���I!�oLS�)37J*u���{��}!�`�(i3!�`�(i3!�`�(i3���w�P���+��o�.o�`��K5�w,��"�����q��l0\4L$ֵ����門�ҋX����Q��C� ��!�`�(i3!�`�(i3!�`�(i3k��j �%��:wJ~��r�=��uy������I �P2<WV��
i�c�rד��L��T7Ê7�E�4'���Xw!�`�(i3!�`�(i3!�`�(i3!�`�(i3 ��ii����1��뜙��L`Q�
_�J�g�J�LQ��wEOJ�uxm�!�oLS�)37J*uc�A�L'�t�Otj{%��ߛ�8���/��}�Ш���my$�N��;� ��b�� л�<Ct�a��\=��
i�c�r�]���,q�7Ê7�E�4'���Xw�j�7��k�-i�9~�,0=]^	�&�e A7YzE�ˇ�h����2�[Q	��
�Q�}#�ҒIs{JE���=���B�NoSƏw0���|��*��<��z��}�0z�cUL��լ[po���̛i���7�v�ԯ��Q[R�7�Mei|�{LZn�+�m�&(|dPSM0.�J�a3mPy���dn����]�!��	Ǹ�y85�&�;���
��#E�>���T�\ �͘�f��p�b�z'hۉ)[텡#����Mei|�B��Vj��m�&(|dP`�,����}];�SS<-S�N;��0�"� ��w� 9_�똣w�ٽv�yq�`0�|(O��"��"�T�>�#�ҒIs{�D������:_�_5:��(�I>�IP�b������:�kR�$fOyQ��������b^��ɮ�� л�G/1avQ�e�b�����,��Z?m��r�գ��(W�{fy}P��B�wo��<�,R�8Ġ��x�6Y�nlH�I<�6�Q=���x��<�6�Q=	I%Mq��`Ҧ�׶!z1��,,ҹ�$�OD��G͘B./�<ĩ�46�;:��/k3gS�yy�ã��&�զ2p�$�W��	]�	���F���X:����*�`��g>~qA��@����M�P�;���=����t��LӰ�+M�ҋX����L$�����/���NM����s�٩�삂��!O@T'���Xw�����U�VA�ڦ�c4G��.���"������O�69:�BF�!���q�%��Ro�����:,:��G��.��M�zp�p+!�`�(i3!�`�(i3�ܒ.���T_�[�S{�o%^�G@�m�񈽢d@ǚ��ظ���K����^W��k����I�!�`�(i3!�`�(i3�Ѳ��aS�!-�+_����1�"`��Ę*��7��S�S�yy����9K��r|Z�%%�5�_Z鎬����=���ޒC>��}Dq�f�B)vظ�u��o��C!T*p�VU��Jp��T���ȓM�Me��d	�A��7j�!󊾵�e�;Pq]g\ ���ǋҠ7�	�ߥ�H�^ /m�6���<�6�Q=���Ң�Q<�6�Q=	I%Mq��`Ҧ�׶!z1��,�У��a�p���L1�%�1��zo%M|�e אN�ʡV�l��� л�G/1avQ�e�b�����,��Z?m��`�������VRj8�@��"�VGN�Ar��$x�y�ˏgԊ���c�.D�#�ҒIs{�>Y��}�:_�_5:��(�I>�IP�b�����LQo������R��H�O��	�d[��K�pHj�4�\��F���77AƐ^�8�tn�+�e��j�3����&Y��V�贅���Ǯ0��]㯟B./�<ĩku��j�,�J�2��s] U���v{:��h��MB��V<��z��}�<ͧ�:|��b+}y[�MQNv�2���!O@T'���Xw�����C�VA�ڦ�c4�5Nleo���_�n�<��z��}�<ͧ�:|��b+}y[|�\m���SLq�N���])���/�Z鎬����Ĺ#{��ž_�Fȼ�Ŷ;���@��O���Z鎬�������(���yf4l!X�t�<�'`ٲ��hN�Qa�T�\ �͘�f��p�b�z'hۉ)[텡#����Mei|�t8�0�=R�U��Y���D��L���Ζ�{Q���A���I��{l�f|��rs�i�Vw�C�-�]|If">�7��	�y^�V]��}��ł�!r�dN�<@Iv�,.9������:5A��p��1����A��:��Q�
_�J�g
�z��+?�����Yr݀�@6���E��~@�k��ϳN'v��(]�(�����
L'���Xw�j�7���1�)�c��,0=]^	�&*��/qRrF�d����M�`|�H]z��l$c��"�
�Ԕ���]�!��	Ǹ�y85���`*uӋ�n�_����Cҷ��e#�ҒIs{�M?rh	�L�vNd�)i�M��5�	��D܂�A%Hy*��(&�L�ϟ��7�4C���6~!ոA2t\��{k�h�+v{��lw	L� �
9CL�x��m,"�J�:S�ٙ���O�Dw
�
�{��_r�e~5�O�%E#P�⒍~��$�x�Wt!�`�(i3J�a$�Y  �VBD�!��"��{�R�ܯ	�J3��Iћ<��!�`�(i3Ǒ�e}5��Ь��z�����ҧ���!�`�(i3:��j�3;R�Zם�³5��&l�����#W�U��ظ�d���!iB��lD�L��&Y��V��^pj�φ��<�6����pIy[�����:Fa�7����Q+��
ņANL��ʡ.>�#�աl�P_�_S:g�RMm�o��'����u��r���2��}��]z=2�4C�[��J��I����~u+�uB;y�� �i�� ^C�ĐHN��R��bP�63Z�t�Fr��j�aq4cn?\ٿ�6�Pfuw�w���*y}ev��ɿ���!�`�(i3���t�T�V�r��}�Q'݀�=�յ[+8��H����Aj��t�35L��$
8��2�ֈe1tSjv��wӨj]h�jsrCm�k��At��D�������,�N��_A�y����Q����.��$��#�_wU|�1����O]��}Dq�f��+��9,(W ���t�1tSjv�!�`�(i3���,�N��_A�y����Q����ݚ�Н�!�`�(i3�{3������=���f.K!�`�(i3��m�~r�D);�OA�uW���%K�ID����k&��At��:5A��pfĉ>99��A0ok��fĉ>99��A0ok��W?�;���z��O���p��!�p,��G��z�q'&�!�?�P�����;�|��[*���I�;��H7�: �.�g3Z�j5�{��p��e;�aT��3G?�d���&����}��6�v'���a00��܀�������!"���	�wT�*,��[��7%^�W+��W��a�si՝�:��j�3;R�Zם�³5��&l�����#W�U��ظ�d���!i����ҧ�.�UH�`A뤭��9f2Pih{#�-eɤ,d��� m�DQ3�z�sis@�����]����n	l��Q;�im��ȍry��	�|���򺜶"���Y6�<���zZT���'/�>!�`�(i3D�c=p���%��:7w�Qt
����+g#>�!�`�(i3�?�Y0�
si�O�����rRV��E���ci�WT�/@���@hG���jw�X���;�줦�ݚ�Н���4tBu6�]���~��4MT2g��H#�"8��!�`�(i3d�hb{;!�`�(i3�F�7��Y�
�cc�V��ݚ�Н�����$G�}�U���)ύ^��R�^Ƒ��f�?ǉ�=:��+���ǔ#s��lxj����R��á�~O��&�C�/��x��&^W(�������$wq�����0��E|�,
�e�~w��R�)d
ӳ�e����kn4@Q�/�!�`�(i3;3�����U젩`#�4>?� �1Zt%��m&<g+b󆤐=��n��y����?�K?SƏw0��|3�o�%,�2��E�\�tP�;,�ttT���-���*��b=��B�'��a�kt`�/>N0Θ��ݚ�Н���9K��r|4�:���m�
��,!Y��j3����:�"���g�Hn7�(�!�`�(i3���P�Ƣ�{��WӠq'&�!&R$/����ݚ�Н�����Gx�6_s/֜ yE֩�&R$/����ݚ�Н����&Z>0���oC��� q��j�J^/���i� ��.�g3Z�j5�{���N-{�
m9�Yt6j�"Hs�Cx�V�x�L���|/��RU��H��<�CH�A1m������eieK!�(MbI;��|B�|��X�?��+�|EYzȧԡ�/$a��F˯�+)�+#c����nS�3�ǻ��d���!i?V��j�c�N�4��@Dx?IJ��a��L�x��5��.�g3ZrZ�0m�\�w�|J����;_��8W�w��fD�W�_����ڝr�F`��*>rc��08�����4C����#��̻�Yi#���!�`�(i3(h�+Z�RL;p�����@�ۻ����4%��0/�'�al��p���K酦z�Gb��P��O����Y��(�
t��Y�{'%s�Ǹ2����E�vwx�k�g��U-�eI?��b��C���/S�)37J*uG(�~ �,���cZ�����o��C!T*�q���U�<�F@"~�@� ��<��z��}�0z�cUL��Jv(K�V��c�4��s���o��x�8���/����\�����A���I��{l�f|��rs�i��s�٭�`�̳��i;��m�S��T�\ ����m0��~�bO\�Rэ�ҋX����7�8����u�c:ɶ��o��C!T*Y�{'%s�Ǹ2����E�vwx�k�g��U-�e��{����w5���ݗ��]����$)@���S��?�FH�$a��ma��bft������y�;���g����0ж�~a��bft��N���m��;���g����0ж�~KԂ��U=��5��L�����;�줦,���<C���O�G��o��s4k�r�j�b#[�o����x�&��'�|�7����s�ݺᣄ#��̳�y�5`P�~�s��hvo���$y̮�K��v �
VWk �0=�b ��"r1��?t7u�`'s^�`}��AyE=�b ��"r�?i���7�|s���q��W�qd�'��n�1��ņ�}h$�ɹ��I���x:����aR�!�`�(i3(T�流����>�SS�]n7A��^⠻rRV�������.�lz\�Q��?s�_{X4x�]�V�����TI���0D�Ub��g��~�4�"4D�/�k�_�|��|�7���@*p?{n��*�LNm�(�V*�u���ƸL��؅��FJ��o�C���j�R�s���-&J�ULnU�x�]�V�����n�l�z��q]4-�k���n��F[�e.VJHn��z�ʨ�lC!�i��}Gz���.��6ǿv�ɢ������=���a��z>�n�S�['Ȑ2��;�Q~���A�U� ���_Y�VN�=��i��}Gz�������vy�|�7���@*p?{n��*�LNm�|��yf{��������K�� ���i7�ܥ��2�/��:M/�CՐ3��F<@�Bcj;�J^��J�Y��h]^"���x�]�V���E�(�� �TYD���`
^8L���o��x�R5�A�yx�]�V���E�(�� �TYD���`
^8L���o���	L]q�x�]�V���E�(�� �TYD��BY��I��O�䓟�&ݏ��A�7�ܥ��2���C�0��(����і�Ʒ��u7btcǹ8ߗ:w��@!~�X�X�]�v��� л�ԭ:h%~k��u�������b,/^/��ux��:S?v!�`�(i3�E����F���8�TP--M�pu�����]��!�`�(i3�d=}b�TY���t�!�`�(i3!�`�(i3%Ah�%4
>��XP��ȆS�%������=�-�o�F[`3*�!!�`�(i3!�`�(i3!�`�(i3�b9���:&�>��s�� �5�v�^*?�z�̒�7�dz�H!�`�(i3!�`�(i3"�,�>E����\�v��_�R�G���Fz�Ͷ��>��9	�F(�Z~}�U��!�`�(i3зq8�Ј)w�<�_N��M��+?�^qk�d	��2Y��kک�)��j)yc�n�.�_�t����ˑ���M��iT1Η)say�s��l>o��|���&l@�[�ݸ�OK����DK7}!�`�(i3���4����4Ieŉh!�`�(i3!�`�(i3%Ah�%4
>��XP���{���r#�LN����p$`�̳��i;v�f7)�!�`�(i3!�`�(i3�b9����4�6�t�!�`�(i3CH�׳�B%