��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���^�F�����b�}�<��S�����h\y�ӹ�+Y$�X5�%y�:�8�����;i�%G���oKp��5�3���=�l���ˊ΃�NA�|Gy�W�6;�E���f9<߄i�XTA�3vv�OW�x"��G���r�z�zʔ�t�A7��myOU�<U�2��qζ��'і��[�w�>\�����	�7�c78�o�N�𔃈�߅�P '[z3��j|��c|`���bo��O�%��ѶYɿO^�O�=-5X��4-; ���^ n2c�瞾����B��?|!�&y2�u|]�g,��|���*�)��}N�;+����'�'�p4�G������	����OR��Ɣ��?�^�<Y��~���`@ke	���+S .��a�5D���Pf[}M9"	�0��j��C�I��e�2v^a���s	��7+��w��[:b���٪�mϾ��H���3�{��H_q㝻�����Rݵ �̡*"��{i=�O���sS��U�^����V�)R'�)�v����Q� p��A���ӺQ�t�,��wR��j<Rl~(��.9")���\��Y�\"^̞��ǲa_>Q۔�<�v$ϣ���U�~kP{N�UZ�P��Ǯ�G�$A��_���]5~�*��b:��nNû�ɤ?���:�<ՠ��S!��Ɋ��&��V�!�Z�2AB�'��1=_y�y�M��4̘Wͼ�>V}���VԄ2w��T���r=恪��[��l�+���\�r�(� �`�p��@�)`���ܮ7g�3�5b���3�;��K�2�lPLνbg���Yi	%oSI�$�a�*<�gb�>k���m��_)-���A��r� ��V��W����#H�:'���ߑ8�T^�K%c~~x��g���l�m�a��x"������ץ�2) F�Ϥ܅@`,�����t�͑ö�w��W_<��bMH��J6+Ϥ�F�>�xx�A=��|b���A�O���brF�� ��@�O��!�"��u�|B�3xK���*.t��o!L���I�oV�~M�~����1�圆�8��7�"Y�ҷ���̞ͯ��a@�b�l��Q&����u��E�����7:2��d�օ�)�O+��;�x�:W"΀��y�I���a~�x�Ѓy�3�f�&[^/l��X�N�@�>��V0q�13��]�_���m��U=�)��� ,�ә<���C�4��'�1XĵeiW�d�4���yNP�����u-],�T���3ǭ8�t\N��t�;��c��VKdbL��Q���{����9W���k�׿e9fSM;�G��ھ��_'9����;%�nfgB�o��C��Bt�����(z�*�~oI�ޙ?N������V.��4��@��uq�9��%F����3��Xy
{X�؃)��J�k>�AϏ�9�$�X�7?-�Mb�z�?\���v��FUܖ�)�%��=b���y���,EJO��u WC����*�l,����:�i�p�ރΥ�TbA2B�ߖ��D/�U��sf/2�*������[h�z�n_n�R�ɺ�trT��׋U�fq��?w7w�ȑ����"�_��%I\��*�[B�2�\ؐ�9�����V�Nw2����WG�QJ��T����G�"U��mܻ���A���_��`�yޗ�'_�7H���qՏ�[��[��&��c��)ה�;	T6P.U�.�=�Hv>6{�y���BwD�~����ff�������(�(	l��h҂�Ư*2�A���V�aqa"E4�n׹�)I��_���@�=ϼ��s:>�M	ϿLg XIbfT�8g��HU�YP��M���E����
*��K&y�}�QEv�SA*Z��f��^p����q����p�eԚ^�qNȣ	�%��Ac��T�Bʃ+Iڵ�S ��
��1���:��YW��\�� @���,1����TŘ�]�"��n<�;P����{�+�����x��"I�OƇ��-�{W\��ez��]J���F��a���KX�W�d�[��敚���1�Ӡu��0�fB�*C+Ik�ݰ�~�����W-��T<�z�e߿�`3����\�cg�U�\5|����|u��/+�?˯��ߘ�sC��;��ŌfطL1�.��i~UV�t��S�}f����?�	�p��O>�X�[�!rzy�QHy�L�PX~�)�h��i�YUCy��ܻd�♲u��8���?@G�s����!�ڵ݀����a%��Q_s�����40k�m�M@bF�T��F�س����$(͵�˷�M������_�?��y�Z]&ᵅo�1P�<F
9�8-�4"��J)J���|�+l~��/��\#�~�v��1L�ȯ�ɳ{>��u�Mm��v�=f%�[BTq'���/d�9�>|D��,g��Arq̢�S9M
VC1;0���O��|M����T���#��n^�K�h��6���4q���&�����0����|��"X:c���G�^K���)֔O�z���P5�g����c:e���~K)����]&m���gq�X��CI"���|6�wc� ݡ����2��DS��A�F�Tu ��3�G��^ST�NA��V��¢C`�fi����4ph#B��]p���V���
��}���:�[���6�h�@��>i�źYD��g���ȄT��ng�Qd��M�h�ǐ�.P*�*<�e?�+ybXt��A�X��&�NG,N���
e�E9��{k�.k��YQ64����+�t�������i�
<+�aH�e>�;UE�� ˄Z�>�48L�yzgQb�j��$Φ���/O���:��+q�LK�Ѥ�E���[�h�[�:h�	z�A5*����Җ�SL�t�����=ad�3d���mM �s�rc�E�kj�<�
��/N����N`ܪanȫ䮻8S��D$��hLH䬶�S���`�����D���%����������q���t�����nT������4kdߌ��{ҕ��fƍ��8n]x�p��by4瀚�	m�>���'�ݓ5�_��������q�#]�N��f���8����2;�q*sɌ�4!SA<D(�30�4�E��lAtđV�L-�)���2)�
����XuASLf_��X�5��\���,�D�|ܵZ�ݕX��Y�AU���s�3ɥ�Z�%��!��҉e��3�\�`�$�]�,"�	���κ��$���c��}�,��]]c���g�ס]� ,�q���Ƿ��t��g���U��7��$� ��bW�Q�"f7����GlT%T�jJD�k��AfL1%}7j�mE�֯�����:6g�X�zb��r��VUqz����<f�R����.�n�m�*�(hv*�(3�\��~�jz�d[�:q��]�j��uo+EAv/H��lva:�F=M[�.���[jsy��!K��L�^���D�,X
�5��tN ���\~$ό��#b&��~`O�Q�L�#䓬�H��ŏ����ή���:!��iG�o��<��T�B~3GM����'�����Va�@�3��	C�q��ioeP��Y���Fh�J���:�ٰâ���.�E����h�{�L�w����9�P M�s{�� O��E��\F��w�x:S����S�F���I�]lT��M������L�Ux�o"��r�匬�9:����|��k��AۿDݑ�*<e~J�W���a��2Bt4-�?�v���I��8ݦn��i`
|"ö$�.o��������Y�V���% ���5D#�����@;�* A^L/%��<L�:�86����A8� ��%� �r��,"ꎵe���~�����Q���9u�`���\�A.+�s�gqa�K�N���_Agh4ۥ���g^S�?#�S��|æ��x������!}b,`�ԉ�K �ѯg�1���)��M�ɦh�z_f?�b}t�B%��!hSXaC��X*L+���L�g�9!fhi�������v�!,����6f=��;'��7Y�Ƣ$6�QC�fI�Vjj�3���?6 �/�I zȔf-��M�Vڠ�g���A�%�އ�
Τ���`��Ut��N�r��N���0�At����>։ŕ��8�*	�7��&��@���ߖO����W�4o��Z ���c�e�pXQ����M#��n�],%B��EįO��/�'[7��c�3��p���]�-C�KA���u>@��yR����9�����^h��T؋�ڶR/O�@M�>�kR�i4�] �_�4U��Z9I�a��'���j��+�n�B��()vQ�(�,Xq����
�o�v�7��{{�,\�5�7z�D7���P,-�zۖ�]�v�y���c	<�� ���_�9+H����n�ܦ{�7���hg�3��L�?=��-�:� �Ѵ��A����G�����leH֙������V����z�y>����t UH�C���Z!<ۣ�7cf1^~Q(�/W�s��Z��Ɓ̯���X����P�+ɽ���	����D����Ehĥ_���񓄲L�޻�Z�H��3���2K�I�@8���_{el�� H�C4p�_�e6����󶽱��ρ~�$	qo�+���h���F�جmuG�H���nY>�eLM_�����@ŮQq��TE��G����ue���N��!���7�²նЀ[�(I����Jʲ��xC�CV�Ҋ�6G�7Է�_V�aG-VBϨ �"�XE	��?����`�K��as��֬��qb������xB�'����R�q#����E�ko	^�M���)
�ȝDp�\�pĦA�n�Fo��m�tJ��̿v���_ŷ���62����V�W�A`�����]R���(�:T� _� ��5FB_l ��	�-Qۢ����k~/���i�
c�:�j�#�dz�T1�LC3�vv�嫨��h�.�膝Hy�O��t7�-̍|ɉ��rn�u�s��#]���jK̂3����ʶ��p��`��h���x"E�;�A�3P�"8H��O��yzO}��l�Y�?�y��,�,h3����ZN�fӹ�3gý���x-L-���6��� ֈz��᣽G�r���Ħ���l���l����EeTc��t/����C#'��gM��4�����QF���6j�rt���B)կ?0�ֻ�����RC��P `t��YШil�m��꫉nn�U �4��p� l��F���MB����߃��i�<-�9`|>�
 >>�,a�=k�횘�� z'�-���v�l����RH>U�yh�MEq�=�]EB<����Fy,�_?�872E�M�;)��pڡj�/��!k�AJ[�e�P�æO�<~�����ŀ�*G��ʏh�<��1���.*f��ꮑ�D�B@�rUM��.�㨥X��>h^
����t�F�(9�k�ѥ���E�*OP(�-�ڭ�=l8=��z�2��	�A	�4�*D�mF��^�A�����q��={\��#���]���NZ�<�<v���M�y���O��~��~Zw���4)?34����Ŷ}���t�`���/�ąo���1f���$_���K�� i�����BFje��6� �T�cfwXlc�H*yuF�)>4߉��1�/�]P��)/?7n��y<����jp��ſݡ��e��`�����=�U�`[�m��[���1q�����=���΍u���k�(�1�!�P��p�(��&�����u��N\h:l=��52����6�̳ D���f�9�'$7J�(C�5��a��g'��iT�Rȣy	�Psr���xG���o0z1t��h���2�M�V�؊슮�;?.��83`�?�{0�.�X꟦�L^T�@ȝ,GΗ�o�@�w9)��v�8wSɏ�on�$����b>� �#�[� J�n��©�ɂN]�T3�����;���V��u�$������{�]��(�y·v��N�c�k*뭬�)��ɉ&bxy�@y��>��4-=�t�71��`Se�˲�I����b#�T�A�����}���X�	ܝ=���$؇o	|w�C�{�q�'�	%Yz��-n�Y0�Yɏ�G?]�ҺQ��O�ΰ� ��Z�m�Y�GT).��tw��{��x_̢'J��ևOT9�j`���Z�}����=��Y-
P�?��0�
ǜx7�)��C����5j�Щ�r�Jv�0�x�[�ת?T��ԙ�[��5g��[��ТTq�J�M ��?�E:�G�9�éR���ĝd2�Uuov��P���^������3�D~&��=Em�Z�#������_sO��%;��_C���6���H��F���q-V{��;HQTy�:��`�(�I����W��"_�06�m|�^ڔ��N"���kTyuĉ�`)�"���/�m�(�Ρ#C8�e���6~�"W�%������٘���;K{��i�v�o���Z��
�y�F�*4R{��a���:���҄�e�:Qh\Z�H�i�����>�v��=�e� a�.��{�=$�Ĥ��e��6��6��)aB��-����<kQ��+a�Gj�|���{��v�"ۍ����Ч���GX9� ���M�wٶ�3�]i��K�:��]�eV�a�+�o�.bB%qj��v&*<bw�^4|�a/!7/�v����v�s�bT"�NH�ÑX��s t�%.�|��ٛ�[~tY�N&j�{A��9?�8�����Fp��Ue҄�G��[�J3�A%��F��ƹV��g�<��ĂEC��'y>���A����T�I>���2{�b�Z�h#��ړ<�+m`��8��J�i�p�PHF�eR�]�{Os��{g�&M�:�^y�[�iG��B�������N:ShB���s����uU�#��&`�A���l�`���Zn'�3�Y�vI� �{'}ќ��@�n���t��q�#3�%�F�jˮfX�dt�rw��ƯkӶ��BR�7vض�}'C��7�+gH�|��zM�	=� �ѤU��u�� �_	wG�����Q�B���:dH�|?��vdĺh�e�v2j���^RZ�G4���M��
�,���k�4�&�
��T(?R5�<�#U��@�Կ�?��H�'e���#��EU�!��3���ٟc'�>C�����1(��r����|�'1qO��*�k*������(,�g�e��I�O���'�)K�NJ�.y�d�Tg5�`�jR>@����C�#��j�����z�c�g�s���P!��,Ź�v�B�/��0�a`�&�� zu��J��
���]p¦�����ɠ�Ȅ��}�ST5�y�t��ظ[�^$;@�1$��?�(�R �Q��4���E�����6������j\uh(k2 V�=��*�ݣ:R��b@Bҕ�oS���u0�T�Ż���
�B-�>��<�^�L���m}�5�(�䶃��.�Ix?����r�G//�[�BEځ�`��g�-���&�)=��g�B҆}}�Q��Ғ�a~�H\.p;Q�{iñj�s��G�.�x<�2PW��[D���� �,(�2�V�#���"��4l���@����w���h1�/S����*[�b�;�iq۔�#��Z���(���d]{|A���Z��b��W�S��y/نv\��v��.��G���\dŐ1�,�2����	�ΦZ[J�J受��!��Px+����b�;�5�OD5ݱG^�-�Z|�ɰ�_z�����8��7]��s���::s�ŨN&0� `)�Đ�Q%��<�<-���v��?�E����jN��L��Y_� �KH����/O���j�Ϯ��	ΌU���8��X���Xi��8����ъg�������2������J�v�<<�P�b��&Ff&^��������oVuZGI��G��1mi{fG8A�(@g۔����k�)e�f�1Y3@d�T���'��ʉ�W�f�� <%�(H�)��C���sIM)�s33��7����O��4+����ƛ��Է�����Q�/���u�,wM��!X�ѿ��lt�|_>60xk�Dȱ�=���(:�Cd�ۉ+���;���\RL�GU�u�u���a�љs}���
�)DK�������̑�QD�?.!8x���I�r;
V�G�f�\f�eh���o?���Q�2 �Ss�f��.Y�u���t��	��m��:kJ��v�]�wl�ʞ5��(]�I5T�����܊Φs�т��eR����Zp8���߫� 9�KU$Yd���ZȎ{�R�n�Eҽ��P�LUF�-���}�祂��1ޯp���&z��村)���=��]�:�d�v*5jC�-�s���so�T�
xTA򞴦T�v��tl4B'�cS�VH�6H^B�V���v��炁�������E�)����]�$�㹪=iO�w� m#���*��h��M3Q�ߧ}��ACx�-أ������!��W"7��-/	x��)�٠'^�]v}D}pP�_���>����іb)�%�[A����>����1���W�L�&J�?%�zI�����w$�g�5H5����@w��Z���g��e���7��H�vy�jU�s��V�m�0�}/)�cR�;�\�����sR�@Y3�����/�>�g�
y�Hw\-
���j[^ɶ�a7D��t%V���)�����{���eҙ�����gڷq�-a�/}a{�2�PgA�Y2a�u7Ʋ���D՜t��!�$��_@$��:t�`Ǡ��u�{�� ���w���t6:.�gei��~�h7ʷF��������-�Go��	k��w���L�T�Z:m���k�3Z9�>>KG���==>7���Å5(��=,��!�q�+*W\nL
B��D�R*�gl4L��D"�Ɲ�/��ʟ�wy�٤�"�;�,5s�f�=�������� ��N�̤՚h�$���U8�r"��7(�k�`ru���/!IxL=�cs���_��
L��B�/�6?���@po���Bi�����o�tͣd�ݠO�/W#�)��e���)���۽SY���*ɿ���#�?p9�01	�S���S�Z����p�C.^�ia-�ݺ�Z9�S�ݍ�s�p�IڥMűzl��Fv����z� �8��e��"���1R��l�S���F6���f6�q^��3* x��9��d�N��-�d�XIZ9�[�"�9c�1���B�-�)}$�Mw�$���7eYZ���`��O��ј���d0��qm`�b�(���:+8��9��"ߖ����n˘\�|���҆����i7� (�j2�y�� ��F�t�yJBP�40��Xz`�T�iV\�c���+�qm���u�M R]A�;��p���J��0������a8�g��;Ej~,�
ʪ�t���`���f(�@����}\�e�4���M]�7"v�M�ۢ�������',��Fq(	b��[��U+����1�c\F�ߔL��]�Z�.��[�	�D�(FL�J��2|GL���u$��GB���y�9�J����$�OƤ���\�<k��=�v���Z�ΠtwR�0�ۏSbiH���8��B�Y��:��`x� 
ٰI�O��+P�r�S����m�\����x���5���/�g������O���Ib^Fİ+��SR��I<�]y�8���
:��^S��.ϳ�%��!��t"o�qe�y�s��46�x��
��H�/6�pL�ި�<Oq��w��i%����j�p	�_M,[�M��"	��c{Q�6C���Z	�2����?� �Z�x�K�-�����ڢ|�K��Omv�G�&[Qb>�w�;��R�C�A����E�Ꙇ��x�d����)�b�b�r&��ԂV��o/��<�U�_�8I��ٵD ��
�_ʜ�\%����dO���R$B�2�uj���ɍ�zP���Y���	Y�̮k,����cD)I �~�O���ڻ�ZIʶ��[ҹ��%�����]{�C/�?��~��!�� ��wX�?�&�u~��ч>H�K��y/��!>�%��cp����~����~�p&E������lzbҬ]�Uq�(/Y�׈��Nh{)1�1�\�L.��'��^�,lS�~&�;$K��t/T�N�6�إ�j�>{��y�]|g]	>�Sz���~6"���[uM#:+wID��MCSit)seF� ֞��$�I�!�=j�-��U,��s�M�q�o��4{�p��y�A���#�`��O2ĐA���u�T�o�Y:e�+�	�?�t�!�#&���=�Q; ����m`����<͘M�v����J�����S��X�-�z�[xIB�J��u�?�Y9��������m<_�x�}4鮡����&�&���O���]�R���M��>W�c��V?���Xdt�B?�n"k�
�ccH4�܎��)�-:����g�";u"Dkl%z��l�o�=�r{��a9$X,�� �_{���}��^���(Scy!��hR����]��#�>9�hq|�T�$�H(�Q}� �� x��k{� ��=�ɶ'���g/�$شO��2i��G�K�~߿V#�[�%�#��f��j�:+��1�Z�����*L�'<�%?=��3�wǿ�Zl'���.�!�U�X6b��=���QLT<�S� �+W���VY�~�2H#���Եm5��K��1J���I����z ��2��I���qjl7$�+�O6���xx��*��Es-��d]�VCF@���W��w,(��2��,n��Ur��A��{N�/�4��YhKi5����ˍ�0�/�L��w�^�����x�N���ޝn��)aZ���t�Z5Lt���S�.���i�k���aɂ�C0d�ࣸ� ��Qt�Rdbu�����x��T��F��0N�DNs�GT���:�h�p/f|�q�|E�F��Cf�!{���L�F�,�+V���1r��H^iK̔-e2$�on>�M���x��s�o8�n�^{	
��ФuA{���0���^�\"��8���n��ƺ-�crl����Y��r����xSs�>�����>}^m�v[��ywco�9���ZЎsZG#�O����G!�p$��6�c�%b)H��q\˷���,��;�i��kX���&�@H�*e2~�t �U~5I�ս�7�-1R):"��o��@��U��@\	K�Wj�"��,^W�@;�|�)���+F���@8����А�<���ZJ>S�3�|�e��}d�9F��Jk�c��2a^��4���@�bD����϶@Vo��`[nu��s��;>��+أ��a�������*~�Wib�ѫx�g��nb�6����)��__�_܉3;�!�(�p���]�rY�t>Mz��-\��q�H���H��M=�x�.@S� �b>	v_|�ű[����&Vȸ��^��ulD��w���8g�o��)
@���X��P͋��O3����(ɷ�NG��jM�������:�M�B G�����S@���u������TS�}�>�F^S)�˭/$�L��Z�o��a��t$k7�>Xu�d6+�ϐi
�H̓v�gnA�j�B��u�r��a®9�����'ݼ��%1�0�3g�&��:?�iQ��(��']�΃]��G6��ηu�`�J�s"v�<��u ���4�I ?eg�	���'��>_kk�x�M~����ۮ`M�@-U#TI� @�4�p>�a ��{"Q��<����<��|�sXk�N��Hj���L^�:/m�΄{�#�(k�ϝ�6�V��IL��OK�`�Y�:�ȓ�q����T�$�p�:y#�}�1c�5ԗ�.Ҵ$_mΫP�������V0�@ur|�=S������b(]0<뿂�t��B4�R��ԟ��̒��B����ӌ��$dm�ߥ���>��:�Wf�����3Ӊ��)����9��=�:%�T��4U�h��g��bkׯؗ�Ƥ�mІ��%���2$R�@-c@���$��� o5��M'�<e-�r�2.f�l 5[lk��~��;�eP�>���_�:
�'2���z��e�>C�d�*�C*`�DN�%����G�{m(��)�$�ż~{����
�WJ'y�}&Z�pq���u��:p~�}��^�G�f�����\y�������!�� 0F��qˁLe�n2>]D %�
t3bN�#߳k�����ʈX$�+�CC�ъ��e�W�T!��i�s@m��4y�� <��)������E�@��g�NBK8!k�#��Q����g�aT)��u�i����eS6�O���&Y�ٝϺ��>_׏M�K�-	2���Q��M�oq�uC���ae�㓬����c���j5��;��$�?��odk}.���Б��Ѻt	[B�t.�l��T
pH�2òo�r<:���D�r����l�i�X7$�ˈk�� �_�4���z��8�C��$Tg~v%���3�=U���@�����0��^��>T}_E���"��h=���Qlq���
�H�:�/I�y�-��:0�&'�c��`�*p	�����BU��H�	��$
�����=t� p��i��ao.���ܷ+���{���D�J��kJE�bZ�2�Х�� V�v�19��*��xo��#��r<��Y�}]�k��#� X�;	n��H�mcV���v=�-sO?0Lr2iEv��,��Ĕ��F�ĕ�U��e����)vҟ�
��Qȟ��o>�FsVG	Z>�F��r�B�:Q�$K��kL�@�t�-|#�{i�-�������U�o�ľ���`8���_9���Lh$��֞kW�'Rl))�}E�sf��vz�<7@e&'�X�6�0��
�9�z�B��Xf65ޗ9f[3�<)���h�����?3TN���ۙ{��=�{p������g�"����%��iP�>|�{(�b�u������JΎ`'�s���������Sp�L��9L|�=��Yt֊���R�^$?*^Y(�J�ǅ�;O��TF��_T�������@Hs}F.��O��6N�i��̦,o�Q�P�����<����>�@X���2�8j]��R��h��
dꠥ�����F�#K��'�9�Ty쀚���;5:��_ݧAA/�B�_�*�[�AG�Jɔ��:X#�-��������fM��:�dѡX����-/=$���*����b�rQ>-p�R�a��]	�{���"f㲭~K�q�D���*x�G�KYv�p"f��`�isSQxG�\@��#���|�h.�m{W�X�M���G�Q�X=M�+MߟBn�a\�K\b�L��� ��h�R����ù�R2����4�̻�3]��\�k��C�!�9��'�������=�g��̌���1�Ɗ Y1_\]26X�k���
4!&��?�t^3Ŵ��I��p(Z�<�����M9�y=s��v,�"��p͑Uj7�0-E�Є�Y�Ǟ��"�c	����ڦ5m�Ӵ�U��1����^N�0O�T����<�'����u	ƫ�`��Sjn�=;�Ǹ��I����E��V�`��Z#
�ɘ ��� [`����y��%?�>#h�]!��3��l���>�_�M^L4���[8�hYUY�9�P���Z���Lu���h��$}�3� �h����NK'pv�!&�G�$/oyqY�M��MY�dS;R�NE$�;UQYf@ݐO���t"�j=c��Z�5*�0��U���+4��[2ĉHְ���V�7���ͧ0̗m�?'��ƫBȊ��<�����&T~iJ�d/�L�����Ƶ������Gԃ ���&N�v^�W��6������t4�M+�-�ʰ��'n�3�/ة��J���K��)�a`PAȑ��o���5��o���tM�5�؄j���{�f�v܄�7jP��Fy\zoM �g��9d�%[IP��RL/�r�vw֥D>�he��00�6'8�8�j|;��7um��ѵ�fɞ�3��BN�;�W�?�ܪ��I1$����6��4^IyU#��U/NH���@�q|�U�gBٛ�pw��IIׇ0� ��I�)>~D�p0\���=�Q�<�ls����r�\��*���#����ل��,�X
���s�M�R���i]��"�q��~T{�ڛ>w�K��q���y�&"���~���"�q-K���C����yt7j+K8i��x��]o��F�?	"	�I��4�~e���d����ܬ�L��uJ�M-�B�;�����o�q<q^��i�go� F$��K����+	��ԫ�eB!'+V���>�{�y��,�����a.�x��v��f�d����&�	�� U�o��rg���g~��LU�1"Ϝ�]�v3�U� 9������7AO����A�JI�¡�ǯ�o�9 p>�]_N:�[q�~��ਚ�j���(�A�Zb.��	Ҳi�k��X��|�2��=|%Zn=܋���Q;a��2C ����e���o2X��˼�X=,A9�Λ�g�_�Y�8¥���hQ�0~�=C8��܆�}� ܍AGBϭɲ�
�
<�w�c��&���-�_��%ﭟ�1�j���-� �_�2��@α׷/br�C�=Z�Ab܃J����l'Q4)P�nV	]t،��i����1+���y�z �?��QF.���
k��c$���� sux�zk�#�XU㥄r��W����ԩ�v��kA�ufn����{8������Q���1��^�V�S4<�r�т�0�խe���A+�� ���q�-ڶ�:��آ�39����&�y��{�$��eJ��H�sc�+\�Q�ds�f:^�XAf�l4i�d
�F�φ�u�
$��S�s,��(�r5�M�7F����P�Ik^�N�s���+�F���2�$��d���MX�rV���>^�Z6ma}�R��V�L7�{�;���*���3��W<��\;�I{�C�W�����L�%���@H�S�&��C �0�3��b�����n'P�A�	�R��-�S����#P�p�C�vz�./������*
�藭nN�6<�k���x%!1�R�^��)�?���QwV���l��J�O�7~�{�#O��x#�#��QX����t��F?��V!E���E�lUv��B�[{wz��u"i�����i�e��v~�P������uS��=�.�:m����v2�f�_>{	��	���<�V���6~aj����XLc�X�2������) ���юF�G�d2����	���#8r�k@N��O��L6h�]����|�5��,�%�*Ð��o��E��\z`�"�h�4�.���~Pumj���ߴP�Q��E�mē������-�Q��0�]�Q��n�H)Ӻ6�
Ü���g�;�����	f��w���C��(�b�33V<��j���4�}ZA�q�B�a,�H\xf!� �(���3�w��4���k$�${�X���,�� R����9��,J[��V��g����|��>P����!�GPE1�}��6��J��5Y��ڋ� 6	5�z8�l�PO�������p�f:���(<W52� V|�SBh\�(C&����h���V���o�MV�XGKg\iE�ح�'�oх�T��C�/�4��bIP��B94ZLʅ�á��C,t�޸��Nʶ�`Y2�4�þ�hfɐ�S�V��Y�����`��p1�;�r2�6�h�*cG�Q�7�҆�%��̹���j����{�ב#�";,l�S��r�d��]�t���1��f��Y�|�l�2�u�Ā�B_Qwhl�4'^]��ŸOUοp擯�aє�Ru	'ZոW�t���T�K�t�>I4�c������C�i�z%T��ȅY!_R07	eRU0#�__���-z*~:G� ����^x��W�d]0�����R����T�۩�IJE]"��P;��]�uo�^9d�U�"���4�j���\]�R�NJY���M%x:�wR��N%�mHEΨ�|��Ap.�M��k�D���5,�9v�a`ũ����7W���B$�,-�t &bi��_'��1O�#��:��&�;=�#��y�&#D��)�Wm�5qJ�L;@�R���`U����F�a�-��䓼E�����j 8Gq�@1�^���9rM�{y{�\fel��_�uN��������A�6z�E��`P=FLF�ch�ms�[����^1�� _,IU&�g=�z���Ϟ���h�c`��ּ��iݰ}o��0���4�5j������IvS������F��Ge�(I�h��p���\�;��trQ�[г��5���2�
����J�ao�vi�1-��T��ѡ��8l:�Z`���*gg�<ն�w�5w�RN\G��V�'a�$����{�X���$�l�At����՘K���48���}�R�#ݖ��*����M�u��d�$�Jly=������?4�t�%h���򁯯�K%w/�%-2��5qɋNذ;{�ց=�<9W_��t��!��SX&����\��[�#�!S��� ���Az��7ه7�qBO?�v�E���lQ`�g���舿H��J�j������P/ڄ#�9�b���kt��VO��N�/A��3ft���!T����ل���d:�UfM먜�b�>�?�=��W��J$�:�פCM:����ݕȃ��7�P�_x�oo@�n�).fđ�Z�V�/��K�`�����m>�Ə��^>h���/���7�~7�Y�,���� ��������[F�:�6�� �yy��l�ȁ�)T��[����{��F�92�f�P��O��µ�$����U@�5.�qr���<���?I���'Ƴ�ۼ�h��?MJ��Dᐵ�<C��x_�;Oe����7��{ه,]�'�lNzoY�6�b�E�4s�$��i���N;��>���c�/��m7�My�Вԋ�G%�L�з��t�۠(P�p��T�s��/�[{6�:)t-b��W߲�Y:�J\�u�{v�]�}ja̯c�ά���S�V�'1����j�y�XK��{/w��*��~�?Sد�����͗�����.K-�8y����� 
7�`0en�D�X�'J;����|�Z���dü�0�ol��ocGc����0�<��[ n�kFgJ�8"���[�$ꖎ����c�`/��E���L�؁���5��Ӈ`3�g���{M}��3��I\5qS�6ؐ��O���xd�L5��J����G-��%�/l[c���Z����,o���6�P�3@����� §ӭ�Z������};�jS�kW�z��F�E>h��I��1-��af鰞k��8[��< �'���:%�̤J�XG�YP�:��	�{���䪟z��� ң�`�"HL��	�m]���AS�)�����Z�U�F2F:U�6#�8���i��+w�\dU�����07o�
ͪ~�c	d=�[�� ^�u�a��o�j���͓�l��	F��l��,|�k�X��:	�_S�=���K�<����8�A�L���)P�8MP?�_�	�aR(�����}�ש3�]�v���s��!' i���2��2�Ŀ>�H����.dS��i?����;�5�;�Dxp��!�|h[=?ޥ V���񲳶���D9$�F9+9,���G�IP���"�T�7r���o�{V�	��, Mo_������W�}�y�8<� ���!B6E	��;�eú��K.C޴^,����p�A�~Ub��1�{k�{`�t���@��|�ck`P����n��^��V�!���8��'d6��x�х.����/�_�������-H�U�ɬ�v�{�]�L�v� ���yIث����Ŭ_@�P�B{q�j�փ�Wi�'Ȍ+s����a�s�� ,iַ���R��F��؁}X�F����,�԰�;y��H%�YP�(��'�#5 V�oV"��J����46k���g;z'��;�pQ�OǞ�d�`���U�:�K
w$�D�XA��������*��(�SD,��^����e�ư�.! �� �y�9��y��%�`�"niذu�!&H���1��@}�XߚhY�`�֝F�`;)�)��U[!�X���߶l���BWm�d��|��K(=˻�hL�����y<���j_sY4(����ATnG�C�)���1tFr��!"��ʷ��]�g�kNx����AɁ<w��z&��CA	ܑ_����J=�$MʃouS~�%�0E�$�$�"йᠹt�3�oe�:T}��}���+�w��{��8�y��Z�SkǳJ�<��va��P﹐�� V�	.���&:�΃�8��P�:	����dR�ќ"#\
lr�5��d�����9�P�H���q��U�?R�h!� ���h�`��|�-huQ���Zʥ0�]�@j���<L��d�@��M�V�C��=�&�A���{��D��Ă����h�(�7ǯ;�o����_c�¼Ї��~2�	��m �D�N,$P�}�Np�#5IR�Y/�4�����՛.��m=Y/�It�T8I�J���ٙx�9O�1;���_.!n-�|Y��AqF��|2�[yQ�Js�'UR�c��;��"�3p���r@�Q����bl�&���J.(Qs�N�#��E��{�P��J�	D ��SG�>�Y�B��#�OQ���['���x.�T��#.O�%&Ò
vH5��$̷�������ʍ4^�UR���x@��e�Q6��-��}�b6�����k���_����
n������&��@��&��S���]�hy�S���W<�����_C���o�h��n`�F(Nݨ��mZ[�4v=l�F�=���		�b���9�lJ( � ~a1�ڣ���iIA�\�����u��a��E ���v0���0��&4���)�bV$<�4�]��S�]��y#�����n��I=��l{�=�xaN9���E���1�7��m�䤕�.L6bvI)�Հ'A��A�>����*���5̕w�1C�F`(45^�<��ғNqg�h��]��)W�'<���`ܭ�e�0>U��N��{
��.ρm��ז��H�@�,k���A������U����l�3��X�5�;Z��9�+���k��7p�Y���+��ldr�
 ��Ԁ�¨�ٕ߁��?�:;0�ږ|�'W�N�Gs;��d.��2CJ�͎1��2�M��f�!_��74�:�p� �U�t��8��|�U#��.��yA��,��/�v���+I��VRUj=��hV�t ؀ZJ�Km�3>(��Z���Sb m̛�!���[~]S�8���%ȟ]�3���p���}'�W��Ai_�s�g`uW;MD��1E�r�.�K����T�Z\m{9��@�+��
���#������d!ys���fÛ'��5a�tǃ-�<�Edi��秝^J�z����k!�b���#I���v�Ԕ��-���l
ۇ/y�K��������,^9X��R&=0� ��g�W��'_�3 �RR���-�w���!>!�a������m�n}���0m{��+�����w�a7@��;nu�/�P�4]�3����XR6�KR���V�/3�h^���|	�M�0fr����<ˬ�4Rv����Ϣ؉�]l�pœ1E���l�P}t����8
���r��E
y796]�����l�3?ؓD�����%G�x�����hOC��ta1��/	�:1\zl���"��;6�������Ϻ��m�H�?b����Ll8.�X�x�H��nι���r�3����A���˥G:���q����_=-�'3��4pqw/)�l\i��;�O�T`�>qz�\[�5=�(y��x�N9*�n�y��!��?���߉���Ue�Cb7jl52����=Ғ�VC�!F�TiKۊ�OE��Vr��~nӄ�k���D	�3�5��/Ӫ�g�7�г�1
���uh���Ϻ����n���"���i�u�y�m����X�H�X�m�Pc�"�A��$�T�A7��#:ȕ\�s����<�o	��I���W`�kc����I�Wq�l�Bl�KU*�����Avx�����TQ*��/��;��>�р�Ӆ�`�4C�?�[T���g���&����;���R�5�A�Sk�a�&k)�w�i��u�Mw���ǌ�%�[��:kr��ώ���������5� $�|[��L	5���<���AB��-e�z��T�:yh�O_Mo��3�y@H� �Ѯ'�0��o����mw{)�|P�U!�T�
�$�C�����%�}8Z�X�W����������N�9G���#�e���M�����7�f�7�,� �MV7�)�~sdj��]�:�&cq��l�95zg_�u�s��,��~~�m�}�TF��}����K��MB7Iߓ�h	֧���>�\�����oJ���������N�{<o�acֳke]�Ο?]4�S�~�VjϹ�e�!f�W��0d�&CU�b��j�[rc�:����`K�D���0�Y��,<�j�c�ܸ���8��m�����e��K'P��񂘼QOF���l&��
��}'�����.b��G`�W�hj�+�)���%V�����3�u%��t���
q=/jN.���=�	!w>���F���E?U�:}?�NN�^F� ְ�ϯ�9��F�̣Yj�x0�>�����	�r�\�� {[`l��MN�J�fx}g��n��w�J�F������>���g�<�m.2;$�X�)e>���K�7�Y���j[]����G��H)ݚ��I6�3�����#�(p��. 1F��_=��U��m