��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�����|"�3��>�U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]�~"ɟ�S��P�jh�I�?g�f&:��r-,^��+o�7\F���r��C>C�݂�N$��/���	�0���'v6�o����Hm��� ��v��x�۔7�D��:�b�#�Bn�am��'��G��҅�>I��4�Ҋn�ڧL4�,3���\.�"�K����u����l�|���j^����;��;��0�Ea�ew2�\��?��n;�|-���g]��~����B��Ճ�����:��M����k��GMG�2�3�NUl��Fj�EB�1~��6NzE�5�pb�Hp�ֲ���#���ƒ�{����7c���:�vq�rY�d�"!Ħ_����ܔ�ߎ�
1���Jm�W�R�?��Xq��Z[�ŀo��c8m�a1���F0XvB�U�@�U�2E$p�����po��z���w�"�SȟL��ə@K;�r5M���
o͇|Ù~;s�+ �:���?.�R�0�޼�d�T2�+aPK���_u�:%�}��ɣ&����B�[aO�d7&'��Y_�jrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�'f�ٵ��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l������ ���yX�ئS��.V&��B֥+��@-�-'͏������l8������t�iZ]XF��������U��֜��3!�`�(i3�:ET֤vKzL͊�q��)�0X��r	�%\*��>cZL�/�gCu(o?C!�`�(i3�:ET֤vKzL͊�q�����$�!h!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��5�Y�w����buߠ��0�z\+T��A@�r$�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3M^�Q(ҏ�^W�U����*qsyN�hΡKCh��(	�G��^�����X=��}DD��;���Ӧ��Gjh�rO-�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��������n�T�?��4��y�-Ղ��hV��6�SԂ}ٴ:!�`�(i3!�`�(i3!�`�(i3!�`�(i3E3�����&Y��V��4�녥p
���$F4���F�J!�`�(i3!�`�(i3!�`�(i3!�`�(i3E3����(I�f�E�ƿ�c �B�dH�7D�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��?��}6���d0J�̛�ĭms)������*��?���-)�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i39�>H��������Q��O�G?X2���Y �67��c��;��\�v�T?�7G|`!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lDr ���K�v�^9�pe�1���l��
$��3R�l��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�
ۼ����F#I�%�[<c�=,�O�G?X2�K��2WIY-�E�f���\�v��_� �u�[؟��)�`U
]�,J��)�[���.�3���j�\�"����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�,�-��L�}�x�6���7|)�`j�.(Wx*�_F�k-�!�`�(i3Y%T��BPe.��xu	�>��l%i�-̇i�d�?�!�`�(i3N�By3��<�]�!����M[��Ǣ&��s���q!�`�(i3��|g�Y�'���Xw���ov��ׄ7-ڍ�qL�\�b�`1���40����x!�`�(i3c��Et�Y�{'%s�Ǹ2���;�¬pX��g��U-�e�,���6+�@ E����!�`�(i3�����
L'���Xw�j�7���5�%]���a(􆿳�ؖ��d�I��-�
�]o��in�m��+�Z����y��.�V�k�J}|��XH�����,>$+W��� j+��@-�-'͏������l8������{y����x��F�U�S���QG�/dH�:2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �����9�+�c<c�=,2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��o�u�/�,��E�1M<���8ss2����p[Y���"�$L$E�͆����~�!U���4��)�Bi�v�V��2*Q=F��&|��~��o/uδ�Q��G�S>���Ol�BW���<o�� �,��D+��bc�n&��<,��	���� �W+`�x�o/f��YX�<:���h�n(���˧�0z�cUL��Jv(K�V��W��_�ړ8���/��P���w��a�e56<���HY ���#�$ݵd���lLB��`���;��|B�#���	I5=��H �C#/<���q�]��`4Ƹ�䴃���%����v��ʡ.>�o����D6�~�ݵ|��*�u�RV��,����>�v�䩲$��߭�?8�)<;0V5���'�ZX^�O��E��	��_JI��_��3�\F�^ܺ�ffJ��IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7�:1��=�6�l�Wߓe`�!��:�r$ɓǃl[�Ƶ��I�q����!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R���/��@���܄��� M�혅vº�w�⽒�rM�e<�N���kb�r!�`�(i3b0��dr����ܓU¯dN�<@Iv��nt=:��:5A��p���W0�]��x@���̢k���F�KD�Vr[/}>5��0�7<(�lb��� л��E�BS�+��U�,�P!6�V���p�+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڲ��y��lDe 4G�1����5����y��lD2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��B�w{v�s�Yls�<Ԍj��_�mS8<�n�ݚ�Н�
̛�]���Wj�$���MC@�����% m���+�t2�-6�=����|2;$�J��7�OT�,ȯ�By�`���	�|��!�`�(i3
̛�]���Օ����@`u:j=��ֽ�d�:5A��pfĉ>99��R�V�"�0�
�:qEp:䩒=]'���%>�rGO�D mWN�Fr��j�:1��=�6�l�WߓR�<�t@@ E����@`u:j�mt�[��������]_��)iƃ�;��|B�#���	��sӮ�}�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���߱QD=t��T�x���b�m�On"WW�ϗ¾IŌL�@
�䪗2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����z�}߯�0�1k�@�����!�`�(i3�l�|���j�ߺ]kԬ�;V��q��po�h0�h����7j)�x����y��E�EnkgR���0?��ܵ�S+J�����iА����H�Kc���- ��5�}�]����8�zƬ���I���d���!i*��?l�ǮD���i�ڿ���DCEF7�����S��ȍry��	w�x�P���E�`JcU!�`�(i3����u��ۦ� ~�p��ݚ�Н��^yE⛀B��+ H!�`�(i3
�V_nu�$�F5k0B�9��n�7�Y��ݫ�Q,P�aw=�"�,�>E���	h��IB��`���o�
P=ܽl 6�+��(����ޙ��E����FWA{I�Z�-"{b��~�Y���(�\w��B���!�`�(i3�l�|���jWɆ&6�\]Yƨ@0�$/���i� ��_������ȍry��	k�k�c7!�`�(i3!�`�(i3Yl���#�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��!�`�(i3��-pө[�!�`�(i3!�`�(i3c��Et��q���U��ݚ�Н�4?s����k!�`�(i3!�`�(i3��|g�Y�'���Xw��}Dq�f�E �W&z_���&#ݟ!�`�(i3�]2�y�Z鎬�������(���	t�����"j���b7|#9��+�t2�,E)�ک�!�`�(i3"�,�>E����-��%M�rs�i�نW0��;�¬pX��g��U-�e oȍ�~�/���i� �B0��O2��p-!]��i۩�s����v^�n��Z��G.�w�ϸ��#|ShI�ˋ��Zt%��m&<>��%��JU�a�(�#��Eo�3�׈PzO�e�n�^��u3v��U�DnK�]_!C6%K�pıs��7��!��}DD����}Dq�f���f�\����U| !�`�(i3;/�"���_�����ݚ�Н�.ӗ�r�(Z+�,�~�7!�`�(i3
�V_nu�$�F5k0B�#2\z���&�3Z�K�!�`�(i3"�,�>E��L/���?T�%��^[�r������z�r{]i!�`�(i3�l�|���jWɆ&6�\]1]�?���(��.�����R�!�`�(i3����X=n/a�τ,�e>%����7V���s�������"�9(�����u��ۦ� ~�p��ݚ�Н��>�@�C5]�꼧5#b|���M
�V_nu�$�F5k0B�X�o|3ԁ���T!�`�(i3"�,�>E��L/���?T�����"�!T؍��R�ٓe����kn�N�Ae�#��� ���)�{� �"!�`�(i3�����5	���]���>����C�Y��j3����(�a��!�`�(i3Y%T��BPe.��xu	�>��l%i�-.���睷!�`�(i3!�`�(i3�E����F7G#+�Ǘ0z�cUL�2�c�L��lC��U�T�\ ���:5A��p�Q9����!�`�(i3!�`�(i3N�By3��<�]�!����M[��Ǣq�\E��0!�`�(i3!�`�(i3�����5	���]���c�A�L'�{&j����6��	�\�HP@�a!�`�(i3$r�t�}i	��D܂�A��o��i�7��k'�w� D�t�ZX`
��⹭�'n�^0o�C~[E[N[\.�|�Q��G�S>�F�1��@�2*Q=F���M��f@�x�OC4��/�#�<6��$)Kx�]�V���x�u�Y�h7�mEox���F=���C{���&�(	�G��^��fO�)�n��
�CӞD�|���P�Q!�`�(i37s�9���o��S8��y�)xʔ���6��	���`y����X �^�m�� �?�@ت��������DzL�Y$�J��;"�,�>E���]�!��	Ǹ�y85��3}�@�7"j���b7*��/qRr#t1.����X�3�D�U�2Y�]^U�*�!��Zo�·:��6�JAԢ�a\��F�dH�%k����1nݾ�����`y����D�U�2Y�~��X�:����8Sk���������fZ鎬����]2i<�L�iI9�o�?�d���&�&�ȫqO8u���t�4��f�i�Q<�>_��X'U���PQ��G�S>L�5c��/���\o�x����ycw��Έ�́E�^��>a_F!���f>x�:	�W+��W�{y����M�V<�';&�C���>~�pS�u�� л��]��`4Ƹ�o�u�/��(s��W���l���� л����eacߦ/�;q
Db%#�'�{b�c��;C�@ڊ�2^��	�Z�kfc��@��v�
H�RtV�^�2��Ȅ&N5�E�E�v;��tr�~Ua�Ns~Q�t�ȇ�J�o��_�Rv�䩲$���dS@Ɵ�oC>��Ӛ��S�J\7r��*�tN1�BJO !�`�(i3�'ž1�|�'����z.��W��!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�.�`��ai�9�^��dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�7<(�lb����?B��#Ɵe�*|�÷�Wе !�`�(i3�$XR�QܛOcOZail������&G!�`�(i3��͝'��ɢ�s�����% m�
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��φ��<�6�&@?Y�#yWs��h�G����,�ǰ��i��W�o�g��G��ȴ.~��n�|�_��Tq�'?�`����a�ۅ<�����B�����;Ly q��j�J^!�`�(i3!�`�(i3��Sk,KXx����y�mZH֫&�z�{d$,���F�cZ��K��2WI�B:�E�h���
�(�s�@e4���F[��W+��W�5w�yC�t��=�˷=�(�Adŀ�<J�Rzh$��{{��0ή��D���e|�e$W�Έ�:r��  � ͷ�	���q��6�Ĳ|4����IhDY�=���6�t� �M�z2p�$�W��	]�	�l��7*�6RRǬv�!�_b���o�u�/
�T^��e�;b6r��Z�X��4tΘĤ�58Z���X
 c�{LY�3T�W	�b����������L�	���+�^��BY�B4��$�[��/� �~�>~�pS�u,��G��z0��-���\�8�E�ńI��)���W�w��fD$0��8Iy�.�C`S�@ys����n5����=�r�������U�8!�`�(i3!�`�(i3!�`�(i3"�,�>E�����k��c	��J�6��ʄA��;��|B'O�d��FiI9�o�?�d���&��n5����=�r��x�9�f��N�D��泵UPal�����_�n��Ĥ
�}+TΘ�� V�E#���Y �6IX���cqY�9�sioo��������>#�(�׮陷fh������bB�o?\�z?Xk�V��	��yAsr�7���X�u��ȋ�=�^�N��ZE��s�m�d�tAgo9��S�!�`�(i3!�`�(i3!�`�(i3!�`�(i3i�|���J�+ H�o��/;��|B'O�d��FiI9�o�?�d���&��n5����=�r��x�9�f��N�D��泵UPal�����_�n��Ĥ
�}+T�F��N���t���ɖ\� ���,ҹ�$�vϸ5EbA���.~0�
n���68;�
4p݅.�g3Z�)V��B�1W���.1	Rv�_�-�$�>ݐ��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcC#/<���q"�M�����Z�H�9 b��T�Q5z����b�3j.�;I)�oRڢ�,��R���'�v�~g��?L׾!���G�~�U�`��}��%%��L���n���q��ݧ��6n��e��'hv[���5���U�ID2��E�A�-�|=�C#/<���q2p�$���\�'��!��h���e%���'l:}��Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcK)�X�Z�
�+C��#�+���?}³nly!f a⣃_B�h���Q��`���;��|B]}�����¿��L��r	F��I�d%�x���� �� eLU����R�;��ݚ�Н�����S���� "5�]!�`�(i3�o�f�Ԝe���b�� �cY�2��Ko��1#2\z���&�3Z�K�-�����t1�,LLM���'yf�?ǉ�=�$�)#��I��H��vY�<��ݚ�Н��!�Ȁ�k)H�=gq���{��W�X+U�"�R!�`�(i3�am.�!�`�(i3y�F_��Jb�[����қDO!�`�(i3���ȍry��	3Lv	̅���8�u?��I��&I���0a�Q�!�`�(i34?s����k!�`�(i3���*[UxG!�`�(i3��zsqG�zM#��m��:��]]t9�?|�i�Y�
P=ܽl.��n��s�X;p`�����c%�ݚ�Н���;�
=�Ww3i�|��SKj�3�H�RtV�^؍��R��I��)���W�w��fD�G-"ұ��<F� �����D�ҏ�6
�+C��#�+���?}��}�Y#&���H�V��h���Q��`���;��|BS}��X��f5a�҉]����ҧd<��2:4~��	�!�`�(i3<�6�Q=�������参1^膴�I��)���W�w��fD�p���C�SS�q!hG������Y�1�R����0�$� ����9 �K��2WIQ17�b�����d���!iO.C�+��uK[FWp�K#J�$
�1d�9���c�}���L��O���6��*w��l� �g�N~}�g)���c�}����T4��$�'��h:���E����<�6�Q=�e��nb�� :�Kn��u������^"�l�+�7#��.`L+�1A]�V)�5s���Z��m/�J���I�U��)���Y;e�iKI/B޾PscX{�X!,{y����i�q,?5q�U`��GeY��H����Qw�c4~Nr_�mS8<�n!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н�{k�h�+]c�)�dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�7<(�lb����?B��#Ɵe�*|�÷�Wе !�`�(i3�$XR�QܛOcOZail������&G!�`�(i3���n�G����|���x�>�+X�M?��y�!�`�(i3�2��}��e�g��)$�{_8�Y��=�}�Vݨ��}Dq�f�՝� s�#���k$ !�`�(i3p�n��W�/�#+*f���]W&!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��׹�� �ѕC?"���>��f�}�	76�&�;��|B���k	���^;�2� (@:��1�
|�g.��g��GԾ�|/a�ñ��<o��8������ a⣃_B�h���Q��`���;��|B��$B���� n2ϒ�ȇ�j����q�\E��0d<��2:�#�5c����Ҫ��8Sk��aG���z���jVѭ@!�`�(i33��0��e��0�U+�qbp@�HN��R��?�d���&�3���L=l��1�R����C����2@P��k����Q��w�п?G����<7u!�`�(i3!�`�(i3!�`�(i3'U���P��\_9ͫ��ʄA��;��|B'O�d��FiI9�o�?�d���&��n5����=�r������`2��'ѧ�Z,α�)IL��	�t�jGԛ>f�� �4�ӷP�Ϧ^c!�6IX���cqY�9�sioo��������>#�(�׮陷fh������bB�o?\�z?Xk�V��	��yAsr�7���X�u��ȋ�=�^�N
�@�<�ľ�L��O��o�a���e��w.�&�H
�DҸJ�v��3�3k���ܼtu�`4��\1�2�?�Z��?L���u���J�F��r�����؊�"�DGMG�2�3�N
;�p?��,"b�\1�N�A!.��{K5~�{5rQ^5�y�o�u�/5Xţ&�	<�tk�Oȑ���Rl�Vn
*����c��;C�@ڊ�2^�}�)����Md���e��9����ݛ�m,���-X��7��C1ݽ�6G�մ���/����'�6�o8:4�I���c�90�Ǘa��xO.C�U��B��-R��l��+X��7��C1ݽ�6G�xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3&�H
�D�h�����0����;q�"��ӌ�r��.J7h�#��3F����Kq��R�=/ ���we��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 zM#��m�.�
9� ���(ٗ.;���JTv���H����o�γ�ha��o���H�RtV�^#�աl�fZ�z9�Y_䈵vض���sˢ.��.�3��H�RtV�^��.J7h�#��3F����Kq��R�=c?5mx�#���ꪆ�l��Pnᜯ}Dq�f�g����Vq���|����Lt�2�tn��뾦�!�`�(i3�����!�`�(i3@�=�{��5%�iq����/���bx/��kOT
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�R��l��+f���U!#���07��6j�"HsS�~�L.�逜��Xw�T� �f&���#��D<V�-�b�+�