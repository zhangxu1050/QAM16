��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>:��cG���Up�Y^����˚;���"J��+��sc��Y6�f$6�5&���z���������`dcR�+��b\�v���D���ղ:h�W��j����='�5Cq����7�r!��:l�6�Fo���_˪��k��LH�]!��0��Rj/��� <0��s8�$h��Bh�*�J}�'�tEs,:l��)+�o }��m����&�X�*��ĵz�`X���<ZR�ڣ�
v��ShAa�{�$`�qC��=?�`�WK~F
�&~�F�br(�g��`S�"\ֈwC��2R��P[<j��i� �L�.�u�T~���GҦ_�&��9rYɛ������05h�]\/�����Z#1�a9支~�؛+7W��m�h�͚5�Ág��I�rǸ��ƕ��׆`_W�g�*���Q�W��ڲ�AF�~%��6"n���r�,�gjY*����Z�y �.9�5t菚���4�5>"ɭ�c��n��Y�8�1��3�<L�&������
����$s(��,�������Wd(cn�w�'�&��xŹC�JP�#-��K�x��QWm����T�pֲ9���M���<�F�jI "���h�M��đ����`w�cڜlp��iA�;�Bxȴ�\���� �	u��f}��b�S	IΨB��}ȗ���9��r%lok*|R��	�}�'�/f�L�n�7��L������UA�/�Sb��#ሡ��.���/�'�Ъ�w�;��!5�Y���f�`� ��°�J�$�N�B��bc&��ǚ�s��#�_; n�F��
q.d�F�sN�/��(6K�i�0�l�O�����,��T�RE�*���Z��7�1:[�L������蠸���?��7($�<3(P?���Q�u���Yno�6�"�Q0aJ��&^�m��C
��S*��g;������~��_T�H$�5�z�q%����koϩg�A�����R|��[�}� ���&'t���	9��n���sT-��y�:�8R���e������3!�@}&\,!�c��-�T��X���-6�B�X/;{w�}�:�y�rUȡbx2�Y�G>�?Q愙)s��U/�&�у������]s���k���f_s9CL��E��)�Wkv^������QTUӜހ�Wf�*|<�~^s�g����&.w�<@%z��e"gӕk�
;T��
��G�4�&j����;��	�����ƺϗ9P�UAVĺ� �x�B�����D�;�E��P8E_���� !�a�Q:����K�/U(�"�
[�PF��]e��j ,s�@-����J�P�R��-򉙓�j&���X���;!��4ůFɀ6�B8 ��P�C��#n5�����n�u9�>?�$��~V��L�lM�ˀDX̗ �X��0�􆘶�UXTT#�@��zﲃR-��1aLvuŨ�}��>_r��yr�D���$����Zn�g���U>��Gg����ZM�w���R���5�흏xH:����K�X��@����y�81��sKI}��#��$�*��G�J��hzg}��,6��p��I�	Z<4��"3otD��R剓T���y�P��M ��ԑ��$Ӳ�=! _�_��\<�\�4�T� �]��
�;��Y����vS�Vx��\D�$nuz�x�^:i�Fm�tD����X�4�咰-Z��hb��!x�P<%�1
����7P�4dM��*���������Qꍤ-r`K?D�'��T,��x��h��|fw�h'�7Hw�T���J�˜`َΔ�j����2 �R�6����}�����9UQ0��n&�Y�q�5�F�HT9�ا�e�p��Y��Bn�ֳ�Flu������';s^��qu��*0���;,=Q��y0h�J��X�[&Γ���]W#�H�;�1�>P�PۧL�ݺ�=J5���̟�:_ʼ�pp)��^z4�]T��B����?��T�>��_Lr��Z���p�{�0b��K��+Z�^^���.���u��>�� +	����Y͍q�~t5�U.
U�~��z�� ?�[�ZΗ�[$I���
�)�,c5�l�v�}��yۗ��||<��KƊ�QK��ǵ���p���diP�_<E���CsU��.s@BǗ"`u�9�Hɗ�(�%E�,���@L��:��J#D�VdW�٨� w�v�ۡ��(۞�P����M�vckH�}�E�]�x��P���ИPth5?��j3�O�� q����~z�z-�~5���\{�t��es����g�J'd��ٳ�Ov�v�,J��JZGY�l���UJ�r���p�f���@�nFT�9e���'�0վ}��v�1���ևD~�۸$>J���@̯�)�ꑽU){w��]4Z
.�I�����.��}_�U�!~B�d+�U^���jeJ�il���pQA�t�:��19>���7IY��f�^l걐oo�J���*y+h��l@�ז]gR�ZGl������� �>'���!#R?�s��`���R\o�W T�h��Z!��Vk��v_=�����ᛯ�	\������F��{g)�*Z�	���2y����r�5x��KQH���A܄��e�vܣ��a�a�Sa�ŭ�@N�R+��K��>^-U@�����	��c�\9ڙ�Fu �z�a��"�K����k&��e�Eo%�#��C;`����Z�8��z�::����̭̅���2��DW"ͩ��Jc�ӫ�p7����<O�"�d�S����������e��e�����K�� p�Y�p6'��dz�PVMx&�&�I��� [}i�6����=��L<�+�L�v�s��h�{`�"&4'��F���p�YhXyw4�P� �׹�"hq�%z�@���t<M���!�q��|c�p��0�;�v��wvj}��1戼�@2zb�&:w�KB�Se�Eq�bׁ����V�R��F�C�a
��v��ηc�y�aѹ��}M���L�#�|��o�T�M���"����8j����3���z������9����:k1���6q�Gh�5��݌%�#	�k�g��.E��Lz �K�	!��Cі
u��<������6}9�����;8I���Q|&�0��~�=�(��j,�ɩ��N�R|�b-����j(��9�ŏލkS?�ęu,&*ఙ`?�Pq8Gpc����'�)�@����1��Bn� h��Nj�c�ׂ�JVo�Iؿii�,cN/{|���\p�àEd�F�H�Y��ɥ?4b�5�G3�Z�6��ΚF�R������:�Kk���� ��٠���Q���,���׺�;:z'���]��P�)�7�Z=}���q����P�<�+�e����ƞ��M�
M��b���2����j���W�*����|T>�[d����x@����}x���|�#�G+��a���b�M!�檁�:f7��麵�����S:�1M��L��mw ��:K(�Aid~SWL�)�G�Ի%�����C�������%dIr��B��*��!,ˢ��8��&2���[5���&�]*�# vQ���%C�z&t-�m�����ŋ&U<�]V�u��k��4�-�Wݼn��x�fۡE��ÿOJ������d��@�^s��Z �?�P�������Q�i�nc0���Q�y����������Fe򤴇%f�Ƶ����8�LoK�OX _�%�,@���	��iwol�m��F�k���g;�5��jz&����}�d��[B oB��(e�\�ǭ��F�D9�o�_�n�M��x$mg��� h�朶 �W����A4�`25��j�c��r�$���@v{��5E��xԧ�sYf�cΦD�R�u��j�|�_�n؜�~��x
�dƺ�"@àcB�W֝$�Ű17ZߦfHJ����}A���U$,ȇA>��]��� %���C�q���x�:$a�T�<ޏj������:O%.��Y�˦-��W����}�p苬��wݝǪ��7Y�r���`�x�1�5.Z�z�����%���'����ޘ��<[�]�!�ࢸI��w,t�ɦ���$g�@<�E߾6�gQ� ��,�U����2���Vz��eӑ��Pʋ�6�{������6e�5� ǻ�b�w
&x�7i�~��\_�cϐ���ҩ��y,iͶ��T�W�����C;ѲK_a�G�U�룘Y���i���`*QO5�*b{Ѽ���W�V�x����3��7M�W�E[�i4Nio�C�o/S[��m��k��N�O���D��� H���Gr�����<�j2� X+��ye����r?ܝ�Y��KCJ�P';�F���vRQ=�(G0��W�����ٞ]{t�cCBQ��ROU���
��R��.w/�q`J;�~�����l���~N��stS>+�&��$ �����OŤ�,�л�����M� �6z�vv��F'�ж����?��F���F�[c;��i�C�c`��C�A��`��$����j�r��b���y���1�R�P��1�z�))l�l��EO��Ӷ��C����F������4
����ó��ݼ��xB����߄���^��?a�(i�ݩ�	�P�O��%e��qU�P�M�|O����n����VBb����PDN�_���;^�����w���p�xkS�A��W%�ш�̥�wٚ�U[(FsD$�o�Ir�����/ұ��
\�6۟2��=���#k�L:�̣��?�8
��J���.���3\P�ǗO�����(��e!wh��R��F��t����7��$�������SD~���%m�h�R��A�F���nB�h>SaV'�Zmt�}�K�ME�̫eccb?�.^B�V���Z�-gЗ����W&��3�}A��	C��Y�@���;��=���������/��,��/�E���H��2F���z��V�<�����3���������k-H�����s(m�L>b<�4��{� (WM�9~ue�9M��+�l�اIw��y4x?��`@��>o�0����j6\g}�ǂ"4�j�+���]#X�&m�^U���E��o�[y�V�hl(,� �5�:��e�zG4k��>��_dfk��0�k�Z�*��8��1@��kkS�Q�Z7�2o��xf��@`	J+-(
�0����$���P(6 ����:�����,w���L+�C�V���!�����P~����E��8�#�&лl@���^su��guW=c@���$�@0����:6�t�k��N�����q�q�Y烙D��n� #3H�]J��3j�rDܿho�>5�k���	���V80f�k����N�pR���	-��.C<0�>��eq�y ��C�<�`<y�'�d�c&`�}l�0�_�Ӟ�f�>ID��;%�9����
�7Q��`�����@9Nms�~k�۴D��Ƣ�����(uQR�?�����$XR~x@4��
:B[�[x���Fw�T2���A�]{/�����ʝ��:L�od�wu��[v�+qoY�� d8N��3����P����R�� �v���G��	
p��a�n�۷�Q5r:_�XK�dQu�o�-:M���ƊOFOFġ�Jx� ��!W���5F?�Z��nYK�W�}�����]���z�$6�D�gƱY�k�=��C~9�a����(�K}�2tNY�:�p�R��Z�Jӭ�+ (L��������e���J5˼)�bJs��5Yz��S Lpl�El��{���(��ɸ����X���m���3N1���;h�i�u�:��̉����q�� o�!�)D�1 �{}�Jme7*�ul R�S�M�32�hw�<3��;2_�E��?"���]{u-��Lǩ�܌��o�~Ep��m��
F �;&������GUq�k��1�-_A��U�H�R.���~�������ݎ�z3��R��8j�H�]�!j��������������Z���H�"��H/��6���d¥	*�L�oQ^w�2o�bm~����F�z���� ��jZ�4Eۺ���e��	�=2NA����	P�xD����Y]
0�������r���2s�����]�����iP�6�������K�#?(��B�2���$�?e@�#[��iWD���1��Ŏ/�S��,YJB{#;d��a�o��uw����R��wz�-TJ�[�IS>����jf �;$Ђ���=���ȅ����>e�~ƽ{Fa)�X�'q�4,��,��z�M�����ݙ'��ృ�����{g,L�t�(�c�I�S�Ǎ�xG��B����̳М�