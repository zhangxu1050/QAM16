��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf^��$�i�g�Wɐ�)
�Ql�Y�+6�iѰ�^���d�u�.�Ye�ZG�$*�f�pM��Y���f<���YB�H6]��^�8�G{��:RjeQ��2
�ƣː��5JLO%/.�)����\�
,��YIw_�aJ�/��]b<Q�	�AVa4+ط֎2�h�\�f�c��^�x�l��w�,���hw���H����.W�f0��G�s�� J�d������Kn��_E;��X��*�M��f50�38�N9Ga_�#��mV�ƭhbD�*�+�Е�Il�ߕ���09-/�p�暌��x&ڠ�	4���N�9D������tI���K�~�P=&0�L��,��FB��������G��K;��Q���q�m*eP	�� ꕝϓ촅J��&:�g,WOn��7[��*������?��@���;�Og��B/��8��9n��$ް'���j��FA7o�6�Fb�km�l��Ѕ.�qͥ�<�^(�#*� ���V&>~�S�ӻ�ɌjC�0}sN�P�SN�<��� Y 4F,a�$�pe�4��U��8��e��|��Y�J�J�	���_:�mQW��=n������<�� -�ϐ�a��Ih��v!}<�jHV�c%��A��(x���)��{�~��k_��`/��;Y݌GD�G��CM�U�����g������H����Eu�A�[%�X7q֫8Hl����F5����X]3ہܸ�W�h}m�����.���;�pŔ�-F���o.1'M�?�hF�߬��5:CGH�b^���A�/���W����9�Y�h(��:�y�펎0��K�'�e-K��\��Աp|.m�_h�pH��,�嵷Y�U(�_5!:��z.�x})?�]��&$V]L⻂�20�V� r�����,�ʲ�L"�L����#V�t�y��T`��Z�z�\�,���:�D�j�	�_�����X�����Ήw��+��-�6��$�����RD}:�{n������=M%;�D�
�H�G���C[�X�C:<%WC�´�A��?W�m��*��8k(��d�!P]��4}�c?`�������;Y��b��u<�ܴ4������Ky��h�<s5�r�ʡ������Ar֬h�蔽xo|��ّ��{����_��lŝܤ�-����DYt�ݧ�AO�.��Rp��C�k��T���{(���;�ӉSP]��b��Ni��Ƌ�ƫ�M��%1�j�װ)ʜH�o�k���$�73P�5�c������UX�f%GB�۵x��x;ҵ`�H���	�vx��/x�jWOfT� JM}W_��p��-�-���5&I��	\D���.Z��,�M�\�*�X�f�@F�͓��G�``�����W,�٥�}�?q
�X��̯N����c��|�:T�B'~۾�~���r���N��A�"�m����`��J,�Nc5n�)sk�� ���]K`�P�L��քv�1��h����&�U����9��էn"ZWHi�3�·�4���y.��ѥ9ץǾ��b�B��[����Q�������ق������OK�/��՞�L��\>B5�w}	:g���{ )1����Q'%τX|�5.����5�N����L���ѽ  ��,)�2�yؤ_xt��3&���%��$�SB.�!O�pZ(���u`UAk�h�A�L2fZ����%�����
~��?��?V�� h����r����ւ*�h}�iB�-X:�Ȉ=�����������_�#�38�gt���D��'ŦŹ��4��_�:\"�KO�����ft�ω�����VK����m�\A�8���P��a�c�)\��j�	:�Gy���p���@!�@���ʾ�7� �XK��q����{���>ے-;���ޡe,����`&Kv��kWP�D�o���s���g��^J,��%�F�#����`R�<��>d��d�������?�F�@;�q3#e_e-�2����W�l�@H+��F��;�8r����z1��(
#7:�#��Ε�9he&V�l�zn���元+�G��]]ߖix�WH����<�U�}$68t)g�-�M��o�I��N;�������ny *����J��[w��z��)�] >�����mW/�QhI>I����yF�� =�ݯK��j
��*��F�4m����k�g��n�u��E�s��D����������c'wӕѨ���Y.%���fu>��
٢�I^J�T�HM�(IT/#�(~��_�W���U�%���8���I�A�]xu������M];�"�X�*�8�\\����P�>pO;+�0��/[�}@sKB٣sԁR)U�6W����e۟��L�{|�I�' ���H��O�B�+	!��_=ycs�}�tLo+���!���~J��U�)O����[C�� $��hjW��sl3��E����w�^��-5��()w�2�SL����3�/���Qñl,Sc'���4g�#���6�� i�-y�Q��7��6Q@��@�)��Rl�����~z3�1L��Ʋ�E��ۍ~5��~b/��m9T��~���ｄDuzݺ7�2��|X/Dd�R��J���c�<O�Z���% 9�`���2��Z0k;��<�M��كm?^`�p�[bx�醯����:z�����n�`j,yi�9�(�Q��C�w`���5�jT����z}2͓���ٸ�e����V�&h�a��D�uef�K����S�{叕(qV:9�Z�-k0G�D�Q��.�>��S[���}5��>Y���Ϸ�!��i^ŃJ�9�@W�p�ʧ*�%$����������pt�cm�iD��I��*ԪHi�3�io�y��16�e�AH��0Ť�W��yÊ|c�u^���-�Tp�Uh��q�VU�Μ�ʮ͡q�0��91x�k�Nltkތ&���~����#��{�@mg�Y�]Υ��^a�b�H8w�k��8�MNģw�1��׾���6�%��ij��S��ِl)��(&�
�6�Cdq��`�J�4`����8��쩱H�O�F=*yE�WDi18Nk2�QTS�ْ��L\F�Cv�&�^v�T��__
�$��.��l����H	��s�L%!*"���P��ʔp�/���z;���㡜��0��2]�&��6e��T����4��q?��uj�
�X!�7ۊ<�-�vj3��c�H}���8�.A_?H�j<�;W�!B��0"�|�6����Ȅ�|L���2���.����`+�x;�Y`�Nr*�
v�����8�!��S�C�rl�����76.m���za�H��*��
i 09�D� �ϓ(7��L\��C2[(k����N�r������h Ym�8�f���;$���B�_*��3�'w�3��=��U�VM&�-C#����<j�(�B��_��>���C�@-k1�F�l�g�-xҗﯫ�o>��]��,�0�P�F̤�� O�g�#�E��0��p"�8U���J�Rk��_�w��r�8g����p	nz�:�Q�\)�P�ӥ�\�>7Z��$LX��yM�/, @H<&^�Z��e�s��ZM�'�����&RG��G<�B�U��wB	}�%���H����j*�A O���K%$�6��j4��v�z���֪�TW�]���@͂��%��@ Y����J�H�<CW�\�O_2`w���}Wr�L�Ј�}��|�C�{\�G5;#c]����)4�TxA@��@��$7�[
�?�ڂ�$0�����æ�we6�s�Z�NR���+����zi�����r��yg�g��j\D���*;��$2�� �|
DJD3pU��o���>|�ˇ���צ�.������"j���Tڥ6�z�Y�E����M�EEc�=��Y'Ƌ�����ai��I��;]\�J{ID�L��p�3���T��5���S�K0m��e"aV��55��[��Mq(V�?F|�M�>���Bd��b�B8)ݻ���'�T`w�>N��-�|��]PK"8������<O�.'�	�{n�yƙ�&)�V������M*��^!9\�gۦ����NF��ʀ�v2dZXi��a�ֱ[�yD�#���_G�7�Nr܆��p3��I^R�w3��?���`����2oh�p�����'%��]{$�>�[4�,Ua��.�O��$�$g?)�cR�������\����g)"�F!��8g���5�<��zj�z����e.��ALo2D��,9y�3Ps�M�����%{�}��I���~��fk�t�b��R$4?t���%��e�Z��Q�P�2�n�n��������<��H�H<+�g�rc�*5�>M[eY9,�m�,�t�L�ҿZi���n�mpH�מ]@����v]��1ң��v��ī"��nXߖ��_��OL	�I�ǁ��vA5�˯q֊����A�� 1�%��$ |�>bH9V���=jR]1���0t�Od�¯��=N�a
=�VT7�>�Z�8����]�b�Эfll3�_�Mtq�������*���-����!�G}�!o�����A��̈��4���!j�%=@"��ǯ�l2=�,xY�y�I�m32��w,�(ե�/la��6�c,����pp�:5�w�H�m*2!n�kR�@t�J�
 � ��?;��1��236���g�e.��oA��]��Y�վ:�P�d�%N	��a0��B]C*�s����_�]�}CȊ(X_N-,J����v��\�|��r��wZ�Q��w@eU�C�`�j�E��Y��Du�ŲH�XQώ:|�E�j���؋z�j'!t�����Y�&���
������w#���O(p�����Y�z�Sjw ɪ@Y���f��D����Z�!C�)�{>٢B$J9,C�k�-��Ze.L�ի�g�]�s�W�0m��P:��]������_)�B9;��M�e���Ǖ�E`&h�
�Ր�ZO>�6,��ClBg���ԝ�9Y�)c��	���7�:�d��D���=j��4Ԑ<�� .-D�+&k�I��a���;;�v�ҟW=��`�]P�gj���|�k-.�A�πIS����X�4��%o�!K�n�T��/�Q{�@�F��#�������ӳ�X���ƶ��k噿6�ɝ���y�������q�����]���	���w�Ʋ5���+�
��M����BR�kz�y!Ջ�"�C��tX����@D�(P�����C*��O����Um���6�bW�Sq"x�9�D	��)#�f�Q�B�Y�[�c�P�yu�[�R+s
���� �������ւ+B1|#��X�+�d0�!'�(þO�E|'vт�B��w*jQ��5p�=M],J��������S�H@ԫ[cd5��(%�9���(�F���!wn��']CI�v]pd�����a�d x��P6tj7��kܐH]�=�C� �Q�+�����@1��V�����l�}�=k�����o̻1����Y�*�x����D)h����2���^�P��[�+C���Qy�E.�ͭp�+�/����|(E���\���	�R鳧g��x��.��K��S9�6�v�IgΤ�n"K�W���A�jK�LZ&��Ó۵Zy�t#]C�Sc(K֍Uf�:�y�����fD
��Am��/ʟ��aN���S�A�2y����+��^2e��L8�����=��g��h��"C��U��?�l��8���m��׿6���x��.��d�
�x�K���A�w�D�x9~5����A<�v��K�p�]6�10��{r�і�	���O���w"�K$��\�����2�����	�����P�z�hP8H]1����o(�)�����l�9��[�1D�BӇמ>�N����Y��eNf��{�s��C�/,�㓩�g*�mI �!4NU��!��&���(�ӭw��/8��%|̼\���	��9Wֵ%���V��.�ހ�[_���Ǳg�y"�!���X/ �����D�d/k�%!�|>.��9̀5���jhKج��/�e`y�f/��o+Cr�'���+[�Ҋ8ۗ'����u����Gze�u��ƫ��GpQ1Ch%Jo�p[�q��n��E�RO�V�����!�w.��5s��2�۫+��<�I��n�AD�Og�_��G�qs'��k��c65��������;	�]�@s�t�|d{���I�TW9��+E��@�!�Q7���g*�"p��tK���	�z��d�(ѻb0I�@1�4]���(P���.�7��'������8�=�Is�g� ����p<!�[8*�ySP�w}-\���#6P̍������uy���W������,��hd��P.ոmkKþK
����7�?�, ���Xy,�1ԯ��S"a[7�.�|�o������+Ĉ��H6�3�u@?��L>��fJ\���ҌI��>ش�.G=�D��A�?.��vDP��Y�S��O�G�G}�-}u�J"�2D$�&[U������-$���Q�|��T��eAg��Q"���K2s	
�<�AR|O�A��`�w�MN�RR�t�W���vo���F�!h�c����L�$lM����������7�x"/��}�D�����]1טrM����.l�w�hg�3�.
����"	'\Ą ȘW�]����䢼 }4ɇ4��pe{� ��I���S"��Ae#U�T�|��-����/h�~���UOq5Wn���y��AiBs�[�W�ߣ����=�����!E!ykW�}���^��(��O6��k� 0_���Q�x��RlA���5�ɍ!��J8��Hq#:���ɰ��" �Ȁ���^y���)��Uc�r���b4́w�����`1:��4�$�X�ǓG�x@�@����(������gd_�gd�%s�U�^XJ�*�����I��k�[y7!�:�����<�c�Ƌؤ"E���]W��p�I�"�x��n�Yy�]�Z)q�#a&D]��O%ᶆ�Y�1}I��݅���jw�6�<��zk��^���8�zκ��G<%ǭ�����S�	9���;��M��lȤs:!jhGF��>5t�Oar�L�a�-����3�YW��)op2�K�캈�5g"
t��D�|��̹�®���#�o
��^j�u�
���#@	�A�+����W�ƱyX��}W�k��x�!����>טr�)��x�1.��=�ڻr�h�e]%����P�����[��/�H���F��]@�����>�jsCi;����W@=S�x�}�.�������=s���s��)��2B�>v"�X8��WA ��y4�X^��O �~ ��2�Q�P�_r�\724ZLT�P<"�z�v�X"���y�+��;���_�#��O�X��Z�8�s���^��#��U���-_Ȭ{�j�m��ڐ_,��]��V|�:�?$"�'�9O�1G�c`���O�>�J���U�$ݕa;7�9s48x�=��DZ#�6���5�*�	<젛��Y����n�]�Ǒ�yZ�
�Mݦ�욑�־S�nQW?ν^|И6ŚLZ�Mo�"�>�В&{瞏��B�y�v�W3�-�k�mO7��W#_ۃ�)�y���z��� ��
���G3"�*�2��WU�,eY�~�Z�����.�����3��;'�0�	V�ж���z�5ʜ@��+I��]�Z[QIWp�����71 �������\��&�D%?V��p�2=� ����QΌ�O
2�Xt�ϸ����x�V (���>k�;�1��x�&����{��֡1�$���r�3��)a$�:+���_�X�,��Adr�,��Uʗm�5;ǣ����իDN�{��=R�2�hw���:Yv�=�� ��ڡ�͇hc̰8�����IK�)R��{�p@�yp[���� B��2򂆎�}���^D�5A���y��&{�ظo/���׬�iy�qy
�5�6�ͣ��"���BU�x\��H�攛�CtW����O������%����۷}������k��ס��]wQ��٧dܱ������4+G�
i��j��b�%�(�Ba�����6�"p#j����zXf@���*��U�e���!=�в�_ުA���*�z��нm	����b��(��*��s�a��AV\��[w�JB�<��[\��IYk)dM`�}u��ʾǱ+vY���n*q����l~���$�WWz��������_!��f+���p0�x<|i[�O�C�WM_x\�{
�Ci��Z90</@���ytsnPD7qy��"�8b��M!J?b�Kc��-������X����}�.ߙ�R���eYy|?p���~���R��:� �D��ȥ�����z�o�I*q*���.�"z��-��_
�:S�>F�V���f잗:7ee����P�#5�?�z�ۄy
p���C��㌯��aU���C	���\@����+$���
bkL-O�����*���⑩�1���z�*߬&yV��o�y�ް�8XߋhP�#5� +��"��AA�9���B�f��n`��c�#��\�ˇ�!��~�.�V�C2��>!�B���{a#�fP�����w��Z���֘m��o!|��m���Z���G�G��PYZ����\ŋR�|�lͶ	<�3g�EX �&��]�Z�A�Z�B���+��?�#q��(e
��x���fﭖc9�&gL��.61�!�,#�$uH�RQ��5�$!�ȟ]��eA��d~l�2���ׅ�X6˿8��Z��P�D��λ83� s�x��d
�ž�.	���]�{3�	3�0c�0�����@����Ϫ�;���� <&���6V�+�H!���2`xE��t��?q����_�?���R_�(}w���Ad��[��N��W�������*=5g��>�'���!���4���n�	�)C�&���\���\!K�'�ŵiڶІ �&��W|���簶rN���O���f��_�h*j����0�	�ٚ��sh@jl�4�j�M0�:z��Sa5����|+ĕMnX��dl�Z-w�ߔw5��z�`����u�������p�Ւ�
�u�`!���W��L8��!����K'YI���KOAE|<>�%OTB����+f%!;-�h��r�"����փH�{$~�ݡ[4�Ǯ:u��-p2��w���>\��g��޾�E@��"̮�f���oS��txB��O��L�ql�D��V]��L����>M?��%ف[qJ�+�\4��r�~��q��r�q:(U��i��Y�.��zzY)���~�gfh)@���u� �r�*��=���s�^��(@
�0`xa�f�cT�!W� 4��7"�鏹c��̀�=���M��C��� �����'[tl�t�޵2er�Ǳto�IJ�7��p�$ȍ��Lcן�~�/�>���[8�a6�mj�������gy�����GIS5Z�*ǥ�����:�\D n���R��� �6�{��vPÉGVg��_��SΜ�à|
Ǚ��.�9�=̘��s��NP#��ۣ��h�vfe$�1F�}�O��pR����iU�cm%�%AFC�O�_�{�a�`�5d���&�8�%�p��}��쭗N�b+�A�ƚ�xc��qpA*l�`�d}���_?7q ]g�� {�3L@I���?y3���!�.~�2ߕ��i^Uz�s�۝M��:d_�X,��U���k���&�aw
�q��ρ�0�z�pK�(KD��=�����Oض�UA��h�3�����LkB�o}$��{��;�]9����ߝmO��3uS]���(���]�b_��4S9��=(��k����/�:�C�L~�Uݴ6EV��8 �������7��̟�C�q������������=��]o�P�<F��d�^��K	�U�4uW�[�\���p ��Ɋ���q*��`�n�O���ھ���&����-�x��m�}h�V �D��,t"�ǦZ��/�L���;~�fΎ�}��Ԯ���|���%sJW	ǅ���hF�]�K�Fb�NG�Q���`H�R+����� ����x�`x�g2;��]����/"i��(n�u����4V����f(J�(�y��$���͏$�V�Xn�ַ<�cw���"5�2G̝�&�?���p?����������"C͔���b�>#6k]`:]6Ԁ��2�_O�B(�UF��V�;F�k�T�D�#�ט����wu���"$G��	j	����A&�+�d�؅{�C�����������]����x�ݦ��H���d����΢B�T�,6p�ؠӁUe�A����v��L�g�9�͜��K�pȮ�K�鯘2�z�]��rju@��,6�Y�K��+���Ez���O�/�R�I����{HO�*
��kT���Y
ni�c�t����"�(�U9��~�R��vԴ.�����:�:�*�N�5k��s/0{]�#�In��B����i�m��ۯ{d��t�5��w1�3��������'0�������Cb
"�V���{��|�>��H�`��y�F�k]�T��h(/Ǜ4T���IVQ]�״��M^{(�9�m}���,�09|���-�,u�ퟚ�hHQ�}7O�k���Z�o��# ���'��iA�ĩafEI`�0{�SY7�l	5�Ū��󈧑�F	�b�"�a��S�q�6�Ǐ�S5$� SnlE�S��2[pp3h�\��h2���8ғ#X���ǳ[��?ã���*`���<��C���MD=G�].�4U�L�)��`�"!�6]Mm7����A����I��^d����_>d�F'+�ѳ���k>[Ovh���Bu~h�t����z�_��&��B�}�V���[o��Ri�U���D�;�'��o��*�C:$�UW�4�:;���X��tG�2JC���0N�����w��yX������	Ɔ�<eqmH*�o�����6>�R���ݤ����g��6|)� ���2&�
ƻml6�Mj���#z6l�*u(�N��be�R��:��c��|m�AI@e�����������#�zD:�Z�oL�k1�,��*������0M�d'f۶��q�L]���D�qk��t%�Ŵ��c��o$`�w6x�;r�^H�=k�g��z����e����X�ڤ�o�Q��E�#k��s�[�O����O���\[���-�rC��!�Zgio��s�=�vnG�ի�e:����F��T%(�����gu���1y������M�)|��� J���
��]�zFwC�O{�T ��Zp�A��%�8'q�i����uo0��p����b��S̓	����/�v�n�ӯ��a�$��t^��G%QI�vu�U��]�޴3N4�#T��-v�o�q�]�A���/}�B�C�ł��c��t�E�T5�#d�u���v�֦��]R5I���>��
+��
&�[�KRn�$%�=�7�� ~�-���=s
�*���ߚ5ۭ�P'��˥d	�q���^4X�䥉Mьa�Δa�HlR'|�]��Rk��2�k�,�ūp'�<�7��C�����e~�q&����SG�?�K��'Ú�M(�!�o�M]�M쨗�ʀZKQǒ"n��g����ڏ���?�wx��?�u�
��6Z]�^*k��kqG�� �U	�]=[�Y�|�_� +���f8	����1��X�V��覛 ?�kײ�����+/�ܹ��iI,}sJ�'Ƌ�\!���ܥ��R��*�q���aB]����"�M���Ϯ)�
z���(S}<� ڌ��`��!���g�-��oϏ���34��Y�v�I%}W���i�Ls�˹��(Je��Aɽ X���!�5=���tdG��U�����&���B��/�a}f����S��.j�L�0�ُ:�%"�#UT��"�X_a�V�8DM��@̽���,��ڛl�j%.���F���^Ž6�>`���Q
F�} ��p����q�U�-v�6J�xz�MS���_=���̈[VO
�Y�IA%3O���m�t�g���zP� ���b�8�b=���U��X��ֵ�7!�D�5|ڽ�ϫ�b��)m�C��Ήr�2�Ļk�ҽ ᪣o1�_�Gr���>܏���m�0n7�y�A7�U�~.<"�$��lB���vx��dܚ��#�5���<��"9l�����mj�aWEU;nw٦O��p��diH�d���կ�fr��B?b�Y->;ih�[�C��vu�W��6�aK�X���#�y�IJ.X�7�T8���u�!�T6]��)2���]Su�^q'N����<��'�����6S&dk�����1�\�17�|�C}w$Qr�Ŭ���xt�W9�&k��쿅���l$I˜-��C*y���� �F��}C�gR�\��6�Aܰ]�W43��mD��?[{�VZ�P���ͱt	R�o��ܗ�%]h��ej��O�`z�� �����V�i�k���i�ў�P����"D���&#�j�A�K7{�7��x�0�x�
[�v�~ �l�-I�S���Y����r}B����5æ�֊�q�m�X�l����04g���q��5:�3�G����֜�;9�r��e֦�[b��\�?��H��'4o�rZW�$_�ĭM�>�.�WÓa�I>��Bu�&�mmJ�"#��ࣝaH�T��p����%2}X��yh�H	CG������ʂ�^UH�k��cl��	����^ fR>��G콇��� �Z(���&E{�1>(��u�xG�Dי��&�&=�gV���si|�j^��^K=G6�����q����ef���=Z�A4�p���W���ة��d3H��i�؀���x���hfcŞ���-�LI=�0ȾA��,���isH�������aYj��O9�u�u�1?) �Q����c���q�$��sd�W�M��#]W���A�`V��91�7j����@�:��Jo��Ρ���D���ъŏ�6�\w��;���O�g��K�C10qJ/ڤ����^�T`Z�ȁ?}��t>��b�_����H�\�~w��G�>!�.j[,+�7F0�ѳ�d�,mm��#ʘ�d���N����f��l�;�.��?��](�n=Vw��K}��`G) a_9^�㓍\����q�%SC�X S
$VzJ�#�Z�Z�������i�%�v�_�a��,^��γ�!�
d��6��n[�FؓC�'a�a�JA�.4mE��VPD���|E��5-_BqZ3�=�ZB.m˖U�u<4~،><W�G���RDvLb[
Z��qZ��N|��6^yJe�	ό6Us�.ҥ�.�B��i]zy?e�W�W!!��>�"ϔ`���dMp�[����1*�!H�����<AE����;�}-j;�����>#,q��j����Վb���������y5�NhS��|��	�Tv���1N��(�&�#�-��2�Z7��Gjc׎T��(Π i,���W� ����S[����^�s�9`�&DU�`5$�&9�7��L�:���u��vRwt���#"Ă���BO�3[���k�2סd��B��s��k�]Ge��_�W(xk?mT��P�T �$����/!��Y5a猏ؠO҄���҆�!ҩ�u��08͘�^k6;���4��^P|{�Ġ�R#���1���~O�T�0��6t*2������؛ߪk��Y����[դw�*q�'�j��1*#���tR0_��fy��P�l�����!'
��f-fRH����������7���9_^B��'�1���/X'YQ�^��Ož��ܺ��������=]`���4aY�]1�ͩ>�n�<4�4�7���	H�N�!�E8�Pw�������E���INz雉,��/�]����YNN<���שϿ�h^���T-bl��B�;�1�㹪]B?7ӿH���~��,����S��l
��K5Ԡj*���*�oE�g���?5B���d�NY3��8��/��}u;G�ae���v:��X�x�NYuVtRS��{�A�C���qX�m��>�b#�9�T��y�y�2���}�2����u��Qw�KDÛGQ��(|�Z%P򎷼K$��5{�.��x��&����	|�I�Ӂu�&��GOށV�(T�O�R���{��!Ο�Ԣ5�Fgv�k+s�/�^��\�d���D��o�~�[�It��1Y��n�}��ʝ�	�ᩍ�+;�(��UWx�$��0Ah/F��}d�*a� ��8W��h��C	��Uz�á!F���-��'��V�݋�k�#4x��	-�m�Mn%D,o��#�9��<P���; �{kw�V$ҳ~�zŹS���@�R#��c�G<��=�P�e�*#�'���{�ۂ��9Z�9������	���r����%�q��*��!�z��п�Jm����K��"i?�y��E`�߫�x�8Y�h�n���hwh�l{�Ҡ�Cf�{%�D������C/>د�曋}��Dd��0TѦ��BX��n��Չ��}�&s���ئ�}KWDM	a�꧵z�T�=���5�s@��j��˷�`��n1�^�'j�2T��r��m�z���>��zl.S�c���x�`�JO<Y��TG^�d�a��/�W���H�6���Y�r?@�1�(�#�*��"n`4��>>��q͡�o��t�yU��}��̧����Yft�k"�T%��@�t��/~b��Ә�(��*��n�K[j󾉙R|�-��m��I�;c�ʛ����3�gh�����^��(�bw��'A:�~.l�UJ������*mA=�s�^�B�����&^�Ԃ�۩5�MM�fL,��\F��`�(��@u ��b�@��r���[5?<B�-����-�����qf���D�FO;�|����׼�C@V�ٙ�xk�j
�uy�X0:Y��2ٷ�un��%�?��E��c���	ߙ;l�2�����.��f��Hs��D�{�^�|<]�G�Х�״���1҄�Z�[*d��
K@�y�lc'��0X`�;���M_U�d���e���+?~}/��lW��*�⧄�(����Wj�	��8Ĥ���g� ^;gx^5�^3�� ��v�=Bs�u�Y���qv����P���֋�_}Z�L��R�A�.�Xd��7=��(�. ��N�b��gx��9�m�hrl��Y��9 ���W���}�ߘ�S*"���KH�U�$e�*���)��!����m�M��ʑ�E��G�բ:����i ��̦G
k��',�w��SN���V�Qo������j�e��9A�9R~�_������q���T�H�bC�T������������9G�z;"����@w�ѠnN_�{t�V(����À$�&1	a����hJ��w�V-݀j�^� Wļ�J��7ٕL)�`� 0����������~�ر��A@e�����,�]��(G����f�d��MC��7RD������ov�1��J�E^�Nkх��E�I~z�+��H�HrW��J���Xr�J]3!^к�_�K��ꄝ+/*'^e��4�/��D5�Du{ ֭����{�3@뷫!`��Ɔ(�5�G��Jeݽ(�x}v�AJ��zYf/�ʙ�6��iI>|?��Cq`E�&�x��t�m�#\ѫ�Ѿ��J��04���Ƭ��2tDI����*1 ���LO�SA������S��6NэhLMrε������_�a^8�K	W
hl�A��G�'7��.�i~.G��+���圁�Bb��nH�;=Z�ͳ�@�Ȼ�����"����g���< \��_N~"���%(g�ٗ��@�ai�շb��]�l'��x�O���n�=F�Kg�,�&�%�Kc��|߼�c�����¥��?m�:���,�T�����&�nL���~Ry\qe�<R�������]�<��J�����qL�vt��&��d�l7�	/�v�g��~	��������n0�t��0�$�f����S�؇�2)�洛����U[&ǆ;y�J1�-��w\����?~m�g��ju���X�c�22��xυ�vW!�����1h�!�w�b�;�M�/�p�,ɓ;B�R|X��8����>���g�'.e#��@GKS~���gH�5U�b���4����ΖHD�$����kt�S��ѷg˗ʇ�ӱ�&`6��m�P|�?�g�yR�6�<wЃ�M���d�1�����yK~����-C�g
�������g(��{��u���MZ㦾������	͑L'���_IX�[ua�Z#7��)/6^O��S;�JL"d�Q��!Y+F� �����X�� �ӥG��W��P�Bd��O���6�҈dx��\�Ǻ��'tǾ�iHL$&�Ry�D�sQ��c���[��ғ���a��V̻��?Ԅ�1p�0�����+��5��	^'(�}�3P�V�����V�@SB8E�6���)u�J� =�.Ⱦ�~�+��3:��Ɖ��y�E�'�����s�O���Yf�]l}�P���`u�Ռ�o�@��{H��br��Z�����|!���g��7�����P�|��r���t�3�҅L4���uM� �g<4O��$������e\�Z<�
&#d�mU,��h<iA����	h���%�|�Lj�ZP#��~�kV|����a�̉�k�)���N�Mժ�q�TKE���G�q���s�Z��>�&܄�=�B�AY���b���v��]ė�MFh�v���Vd#g_�k_��*zF/x{=O�.�s�2[�B��{=�ǖϰi�V x�o��dWO��bx2�lb�����?GX;�]աlQ�JfFn���9�;�2��Oq��R����ގl�RR�ڌ�B�_]Ҿ�Tq���_~�8(M�Q�Q�%NI[LfQ{�J1Yf���d�A$8<�^�����_�!#q�hN۰��#F���� ��r3c�Q�މ��)�*��t.g����աN��	���?ᓟ��f�ޡ9��@���w=��@)�q��Y���P �8������<��`����D��-boa��P��2��<��� �rH<��D���J�/�1��J7J���y���$_03E�nIHp�o���[��8xκՖ{����g6g+�e�@�<So�[��0���	?`��s�j�K�*&Q^�#��iv����Û�h�ӈ)��Y�/:��l
�N�(�uN���zˡ��}�K^�F[��%���|������:W��w�ڔ�°i��ޯP�<kX����f�B��^2�̞�����H2�T���4��)I`��K����5Ih߄S_�G�
��4�*�e��D9#%�v�e=bP�(�$V���'sP���"�bR�ʇ�?�9��lT��BYZ����p�:1�$ߝ�������&�:q���s9�^���>�$�.��$	�u3��cb0��Ne?n���5��{Ӥn �nL�V#M��G����A��fc����c'՚���Y���"j�'�+�,��m��o�W���&�x/&6��Ē�؂(��S�#&ܺ_�V���j_0c�P|��>�^��HY^ٹE���Ґ����P�&��*"�������r�, ���z��A(��P�:\D	$��/�"w�"���P!�0�t��]��TI�oOxd/�v�y{��$�9m��6r
� !�;�X����R���p}X7����=�� �Z�����1���,t��|څ�C	�VA���$s�^D(	�d��7����cq0��X���@�z0A��r�)���V��:bn��?%2�z�tj��Uioۙ�6�%硙&O���5%���s�P~@��ݔF���1HepŢ�6�2(mg@l����FM7��,��	'{n�i��c��=�zzo!��:{ 8�������(d�Nd)%��r�q?�0��;�Ǵ��\G�BC�9����8��2y΢��PU�m��ք<�?M��O仍f�L��΁��ä�\�C+�9���ҥ�һ} |g�;x��V"Ng�!�P�p�ØH�>Q���m4`U��IuR��I��As�d���Ck�<.��?с�@�����%��:r�.(u�谥|o�>�-�h4�]�eЋH�&�����U�ViG�[+M��d���1�BPO����)��0���͝Qhn����jIJ�͓L��#nB)c��.���L�@6�k�Q��w%ҹU��	���T|u�HY�p"��lڀ�sh�D,A_��4`H��ld��%��zQ��
� v���Ffi ݫJ$IN�$U t�~�m�/���;03H���,εq�5�Ig}�3flM�Z�O��Q��W �	�����8�0'�-�۠N� �����}7��]���
����q^�+����ߏ�F'
Q1i9��~=�Ks�^�ۊ�XW��+Z�о��W���9(Ocl�2�����o�g���I2�c9����P��[*�\�:&]�* /�������dp!D
cc��=���Ǹ?h�v�lX�cx�x+�o��Td�BI��r ��ۭda�I[�� ([,C�XK�G����ص�{td��c n��5L���j��&��ئ���y�]�B��+��Ӽ����*����C)�
a������S�^L�ko:�?s�S\�X�?�V��d��P^�b��J�vCI%���|,��`�I��–s���Ny���l+�ӗT��V��NM��7 �}�D'�H���˦�w������U�M�>}h�	j�JR0V8B�'J`�����JI���gL����PR��߂/b<f�ihǶ\��� y�f du�8�����_�����*�����P��NS1��Y��^��x�I�#�4���{��(��-NJ����מ��⟹�o�������$1�
ĵf�6�:�E��c
��>�`P�	U�T�[((��������&���ʹK[�Bo����;s�$��:Z�߹�	7��<�1h3I�]���P�J䣢,�v���Rk}��hn\�$ꉗ�%��$��|�'��L����F+ǌ�Pw�g�vөT> G� z��73&X�Ň��.�P� R^�@��d�io92�)��� ���Г�����-�p�q���u�:1#��MRCy��Σ$��-m��!C���yD�!G���B�ê��� �@Y�����U��$�@�fV8cw��ϷfC��~dyt];�@�Q����PJD`���MXm�8%e�V��RX�
�tӧ����a����Z�V#��_"��3�z���5P(���\|%�S��~�H�l~�3�q�\���d��s�cAXm~�w\��^�nx��,��1nGk��$�-���5���v5���ܟ�2�Cb�"�j�!+�;�����{vl5�3A���I�g��F{�O2��(,�����-�]�ѱ'��j]�H0x�ذG��(��l
�O���D��Ǧ�7�c�<_��K �[8w��&�&��RЪ��-�?,��I����+6��;�w�Ս�V��F��+W!����W�b�1gXx�C�o���vJ/���Q����}!=��Z�nR�/��?��Y(ޯ�}�]7��bE`�f�0�u��7^���?��l��fD@�oC��jg*��K�\4;���S���\R�������u\�R���Xs3������b��Gխ�ݛ���/�Ɔ����N��n�l,c�e̚[>Iu�Mh��s�B����?Y�N�Z�|6�.�jX��J��l'ŝ�UmS^(����Z��i9v n�ޏ���hG�gG�ͷ!�����x
���)�����n_ZU���4LV�bIn��N 0��#��4Y�O�O�:���=t���p����E��������.h�����gV7}Xk ���A��'�tgϿ"�a�S�����-�K��c��,�{����.��R�="��ҕ����3*&�%�����F]Pv�_���+Ht������n�w��]�>U��A^�
��+�v�P-zv�A!3D]�6�X�}���n�O��h�	϶8z3*�?�LMj>���>�6@~�Ϙ� ��3�CݭT��)-K7���A�g}����UM;7(C�w���AO	<Z���,?�R>��(���Q-�#�q8����cf�O�_���0Ҋ؝�B�`"M{r���p#9H%) ��J�t�ݚ�cy��ß3�J	�6j|�nE�[1UT�W��@4A���a�e��,�Y����KA~1V���E�*,���ƈk�+YҌy���j��j;�|��i�\��Y�h0k��|�~�,���'7�IVN�>d��v�W�r����0����:��|y��iC'N��]C�EXqY���h�m�k~�K ���`��5,����s��7R��z5}��^a���gȫ ��T&�9�����;1>kʉOqlï\��Z��p�2q��xeL��7Y�4яރ�Ih��p�/���C ����[����iv*	��E�G�m'k�� �hW[��^�'�׷�T�06Rޚ2L�q)N
����F���pG��ub�_Ƽ �B٣�t4?�S̂U¡�K�m5��.�	��)}��=l�F�1k�?��c�E��S�N4\B&�n�� ���"ђw��$��4;�'���(�SeG���ح���2-WW\���|k��i9{�G��c%�Ѐy�I�9!ò.Ȁ���d�&+�뇶�3�gf�#m���0��4Ɩ����`C����6o��l���b�"�V����L�H����-H=r2_����k 9s�-��`M��԰LN>4T�E�$����R��-[�9Z�E(��jt'!s8H_,	hNb����x�U����!��u;�ĩ�A c��F�Z�m����?x>I��T��4c�f���]���C[U�Ľ���Man�fetm����Ã�<��k-���|N�\�������n ���3��� g��1XpC��������[3���7��_F��[��>s�v?�=�ry��ݾZ�eJS	�a�/��>`[U�\�8�S�NZT��=�/1���ww������N��4��3<�B��\U���MN�.���H�@�g����Q��ǥ5Ҳ�E�Ӭ�OqG��"ԃ*�9�P��kSH7��惣:�_�y;dc���k��N�,Z4�:���c|X5k �_��(|׻��U~�J�E�����}G	C���Ƭ�E�d��jޑ�ǁ�E�צњiܔ��W\oD߂6���W?'$+���|�YE�����V�J���D��O%�]�M�壾�<R�>��(����R����뻩
�%M��B��Ja��D�lM,�ݽ����d�V��BN�������z(+������a�N���u#��*�;��wO�Um8@�V�a|����"U ���w��	Y�U�'�5,6���G���2)���v�ƏL�
i��J=�x�l�����|.�x�)�Ш!J���V|�8��MF���[X����B��\;�ɏѐ���n����Q ct�Վ�|�]c��I1�֡Ӓ����xMp�uR��Em��s���(��5K�c�3��+ji�ńUvȔ�d� �!�:�*�ڴ��/U��A��2mu�b�����+�D��IR��z|�_�l~ۏs�@|�&2�gt.��n�NsX��[K5Ǆ�nx�!|���:�n���Q2�h�7.�Y�ꌞ�Rʝ'։����y� ��n@���WA�+5�����m^iڕ�X�,�^g�MEqx7O @��{���B�)�3�Z;�Ѷ��?WM���l8t�tl
�����kTyLW��lV��쇐�����3R�p�Xd��_ފ-�I ���۴FZz���e`}�ޠ|���������.:�l��A��~4�J��4��
-f()�kQ�Q�����mY(>�n!��9c��[;��e&Q�F��1��Gj"m��xp�~��cqz�7��4>���(E=��]_�w�m����t� t�^6���c��HV�~8��w�fX���^f}���$�qѿ���)�e�	2���En�&�wǴ>b�a��[�����걣����6m��qqf��LU$U6��U�6�X@j��`%ՠ$'��"NGe�$�*�+#�����n����jWbW������I�������J�WD�j[�T�"#�
t��nJ�V��/�$���F���|�w����1�NE���:
�mO�f�$��U#�/>�@��5�S�)��CF��{�ܤ�]�G
�{!|�c-X��R�KL�� �q�9�����
,�T��Üe����mƤ��������@�>$���..�Ԙ�3��?���H����7�24=+�^t�R��>� 1w��Y&��K���fNl�|�������G�ai�DJ�4�������2�&�".�
O��f�����:�#P���:�n�ʏ���O��Wl胱oW
��๹C��O� w��˙��O�U���/�y�X��|r'0]��f;aT�8,Z�׎����(:$a��7�hM"*���~�p��η�7۔a��"w��5��m�ʚ���L �����4��%�Q��N�����s�64F�]�����D���y�
| �Y�Z/��	(��-�n�q�	���zލ��	����#lv
�Q~��s<���C��H�<�z�2���jː����.OAtq��'�Ү���,�{���Ďl[�������L�ZB���־S�^�h]:�,V��Ԇ^���%hk�����=��x�Ðl�~���rd���1�D ��uo!��~�t�qR������/�C��\ivuǸJq�yh3� �&\����$`�2��y��5�Z��G���w�8�Kg��:s}���q�S�vqD���l��/�5b�V�C��9y���i�R����s&�s�����~⟨X�ϡ�Ӂ�)y����{h��6_'�,��/��|.Ң�L�;�h(D>Y�r�])<�)����5��0�|��V���D�����]@��5ů���Mu}KϵH����9~W�5j�h�f)Pcג�B��J{;�k��+�JF��(q�J$Bndc����a�x�fl��#9A��/׍�p�7M�U2UY#jł���V.�Z|J!��-���b��}xn��t"�
�|�Kg~?��[����k.��Rq��ԑ^�.����c��#�����
��to�B���)"���4��Ŕ�%�8�6G^�b5�A��?(Bgm���S�z%���
���$s�-w� a9V�$T�a�>B紻��ځ�7��خ�yE
�1�ܼyA�oi��c
�B�)���,S���<��{���C�'lV��!������/�ӗ�:���(Xw�O�Ĝ�������k��|�n����Ǣ�f8W'w��=3C̖����a$b����3��w��&��V5l�����l#`2l���.%�!�c���};�{X�[s��ms\��Rwx�Z%�Q�ګEn?J�9�vՐ���ꦐ�J���_2�d�#�(%���m/O"�>ū/�ٕ~�\�	��b<��C�z'���ͽ²������������[���G�ݱ�T�{G���]ncO�F�l�@�S�k��+}��#x�_g��D�����m
�P���'�Co���6VV�x�;
H���IA�3�	����{�C9J���r�����88ν���Y�i�����_��Z�|$Y�Ӏ ~tl}1S�ҿ������"<23�ו���M\0k����΍G�#Ô��`h���/��+&o5��q�z|;�0)���B0��� W��~`.�� g�<�[��l}	�6#���-�O:��^�Uk;VԮ�����7�uM6�Nt��"	7~hQ4��Hl�3MǢ�}�^��H�6���Á'�P�ѳT���xb�7�<@�*I�v� -�Qk���0�&єVҾd�Ui�|�$�l�,�8q��u�p=�ofF,w�z�?��K��t�R�ě�!�mƔϜ5��7�L꥝t�_&s�Ϛ��������:�Wi����Kw��D�k�@n�Fbio5�� ~���EI���FO��y��X��*��^��͕=��8D��2u�Ͻ>df�Q�꥜�b�ubz$����7�\p֚����b�U���".J]���45�`X6�� ��ӳ�ע�4u���q�h�Rqwv���ܔ����h��ˁfK�b L���Jߣ
`��Ծ�TG�e�WK����~2�k����낪�3_W��}%�Ho����T*'�3 �͋>������7��(�):��N�
g�Æ�g�����c§H�;�y�+o��z� IL�Z���r`3N��Π���2M�����NynD����lr�WD�y!ydA���Zv��B_���$fDx;W��|mD��:�R�W
��Քn�ȑ�ʇ@���[E$ϰѴ�o�u��2�����d�?�l��k�{Ϥx����i=}��<(�������{�ȶq��H9 ��-�,Mt�p�p$�yĜ����D�^�����~m��nu�x�@�3��'�y�WnI��|�E1��p���<��m��#����t����.��lh�!��� �h;mQN�������`f�nG��2���F��/����S�H�kJ�J�P��i=N����r�ٷ��BBk��/�6�[�4x=K,)�s�ވ��l��g�5������q���ݿ� ���V����H�1}����G���ƥ޲��Z݂)��D��v���"�@��WҞ�u�ħ�=��L�.��%nn�bЧ�?Z�^cSّ��x�6���>�̩jHKB<}nC���_�rM�x�	��)4�Ԋ5�>��_�\��L��m)��b����a�6T��ϗ	w��/J�t�Ѓr�h[��rm�kv��>��(�hgnx�>�*R�7��-�Ѡ�>oB��ڈ�Ap��Ղ��Z�E��dG��[�l�>�nO�M��u�[٣�H���0�.;ۛ�@:��}`�-k�����!�������~���@R�GSc�Q!��5c;�D�GJ$^����7�X1�Csj��x�Q�x��(��s7b���d�m��>���1�Aҏ�D���y�{1�.����i��ǚ�~�qӸ&y�_G�^���F��"�����#�L�ߚ���}�����W���7�O�n��HJt�EȄ%]z��B����P�[I�My�oA^cO������G��9g�p�î�����v�����)�M�à���P������C� ��T�Lv+  Z�ܿK`�*�0�9X(��0t�u�o�d��7w0����w?#����Ԍ�/���aO����H���D�XKRя,�Pq"��d󣅡4��{Ij���Z���k�J��Ǵ�^��ޘǙV��1���ƄI� 
.�	�y�0ITo�H��UҠ�Rb'?�]Q�ΝW���o�'D�������5g�0>�����������ZbY�,����ճ�qƯ��'03�i�\��J|ߡ��L����g�I+,lqV�6z@�z��9�nH�Y�;֫ �x��9����`�;U����7�c�*��wlD��*���\� S�^[�d�!B2Q���D�� �Ɯܙ�49����z�=�+�����NvǨ���;�|���{�և���ج����(��Sj���?X}� 9�N$����B�	!9Y{��C�'Ս�.�,�"�v�i�%yB_�%��<��0����6�!b�]�"�%�VCF���!.4��y�1�=s!��Y��#���Ɖ{;�u�й��,�%!]M�`Ї����X��y��3omr�X��ɰ5���d��zӵ���w�~�t�$F����VT�[&�x���J
�;A�ߍH\JL{���X������x�q���CY?$=q��JQ>��,���Z��ڙ?�:�q����=Iٯ�{N����2�-X�)�*�+���J��.<?"��h���u!f�8鐈pz>8�P�̒Nr���z�JX�#�2o����E���7$��^�m&/12/�5=+!�Z�)T&����Y8�jΞ:�jd���9DI��-wD+��EI0���(6]��%�Jl5���ܟ���y�<���li��^��O[>�mXFO�󦎮.�T>M�2�g��Y��g��R)�Lp=���n1���������~F\�h���A�ɩ��cG��r��Pyp�����{Mx~�f 3Ӫ��I��똫�Q	5�����.�9���8L�>o�#��΂ ��,��*��J�0��Aܲ�P�{���R�xK��f9�������β��
F�e��K�#E���2�[#"juqnE�m����0�
!R@�h���6�/)" L���L�d[��[�!i�5 b�-0�,�z��	t�2���<1�_~pD,���d}��k�eVJ�0s� ���[�\X�>x�	�W�C�H�˛x��0){�P��J��|_�J3�Ķ+�U����#`��@r��9�4����ڹ �?W��F��xb�䲅�?�b>�m�b*��=��t-3�ģ�ѩ�Y�������0�5T�ce��s���p'�$�k����� �E��.�]��`�'�� l�x8�a�.���Pl��i���7H*�D��rF�#H���q7��?h�EgK���Ӷa'�cTSZ�Vc|�MU�l��p��i�˽��exX��.ț�ԅ�k{X˥o_c�W��3�W4�>eJ�ӛ�xe^�=:�67Q8�!:MLT��e i7흍6���t,�V�y�T��y���؈iS�B��_R���)w�V��
���F�/\v�}$I7��Ѽ�A� [��t���b	��E��:�KoE��bb�i�N��ڍGX4z�h�<��i7���ӗ�@�����H��]j\(���(�o	ə�T���Nl��3�w�xB�l�V(������h�#c��k�Lp�1h.����f���{p|�a�|ӊ+o�h�𘲄z��L�5m*�P�|�l|�K�2"�ĸ�3�"� ���ԫB�΄+؀z��?d��#��0�:$� ku/��@�Q���La����[�N�j�B=ڝ�kQv���p��M�9ќ���\B'���LJ(��}S�EQ��RX����B���_��g���ZV�m�z�cv�̬h�(������>G���+�^��TAGK?M����G�~lǻ�\&^�{�$_ɥ��!0�R��?6�;d-6�ģ������B��]���c?�H�"�hJ���\�_V