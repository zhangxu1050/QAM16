��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�A�O�c9b��2���j�:��HA��?�\/��q�k��#W_�0����J杦�&���£mj��̟鬶�Pf�s5��q�Җh.�k�/��HJGS!]$�y�}�t+��`���������ʣ��d=vP�I˖����T@����)�SV�������Qʀ�W. �g�t*噦�"T�q��+/��l���
��K����dg���Y؂������w�+��|�0��A'�E��Rū�|��{	�U�8^j6��1>Os�)�#	�=j�a]Ϫ�3�1 ��;���P5�I~���������'+(b�s����g����Y�%��nM��0�o2l��_�4YT���2�)̆N-e�S�"��i�M��>�Ŀ(YӻcD8!A��_��<{�TBP��V��0��$�2Ud�z9��b<�h���7S�޴2�m��|;� �Q@R<����Q<�H�˪�r������mD23�LC�Wz</�%�nuB�x`�3u�����n�CkBzi�n��rxi�!^�Ha�5-���잧d"�3:�U[O���]�@o$�'M�+�%��Hw�m
Ƕ��{�T��x�e��+�-[ix庹��x[�'�3��v�}���F|�Xձ�v��v���¯��u�h	p�'�VkH�m�0�<L����q*��Nd��Nٚ;\�����Z�ī}?������Q1T��17��']מ���X,�P��oA�QP܉S���rϖ���ƵQ�#PL�,��qX�W�FT*Y8��?8X��R�+�I�rVA-x�p�|���3�8�pW%��,���������:�@������(��G+W�%_�˦��!�cr&I�#���WMЀ�����R��5pIy��._�C
�p���c���J{`]�=�YJ�F#��ɶ)��\���]a��YtqEc�
���)���$j���O�v^�d��:��OU��P��9�A��AID!m��_5/j'�"��\�K�2�Yz^K��D>0�8�T �6���K«���iB�甊8 �P�o�lt��f� l�4/��p�i�j�a"@<������W �������s��4#��hH�a��z;m0�DWU�W�Xٯ%�ޕ�� 4x���ƃ�.������������!�<2{����*Ƭ>��9�R��
x�XU��-"У�,�m��&�#/��`3�S���ni���uV�Yt�ʢL���d�Sd<4c4�H��A����1�m���ҽ;�x�7]�{�ut	�����C<x��D�⢫A�gJQ�L?�0�B�cc��61��'������q��z�DƄ'���
EL��𤍡F�v��L:���@��y�Ep��H/�*�A��r�,�$V�L��Im��x��}��4չK9��ؠq�A�&5-���`jD��J���2��e��}���`��W�: 򥋀�g��:	������֐DpW��>a�L/
��K���Z
|��(��k>�s�g��D�?�,�O(��d��C6����E��
�� ���ζ�W{������ԝV���!���U!�� Yߕ`ոX������擒��h`� ���c`M���%�y�^Ƿ�?A}:}��`9cH)�<�P8���s�E}1,D��QQ���Oy��	*%�R�z͂Ӆr�p���@�x���͑e���M�=Á')�9�U���C�K�p9i�p�V�嵐FL��(�n��#�}�l!���IJ��d����"��K�4b68p#@�w�E�=WԀN@ŝ�/�,��H�":����a�&_q��f�	,df�V���j�[�`�´�f�υ�`U6o��uu5.�]��R��L�+����9�"=��t�*�[w���j�e�8>���ݚ�x�^�.�\W�J�g�	��;USy�`4mm_yy)[z�� K�#S�K8�����2v.g��ǎM��Ȋd���1�*P���[��@�TH�ei� ,K�M�{���w��	{N%v���gH�]E�҃t�_�0�RŶtM���߾�q�+��%�2�����-���V�o��oP���t�*����pxW!ֻ&�=��&L�����?r˶������Q��k:��\Et�_.y'u`lk�T����t�X$���ɟ
綨�-�V4R��bh	�5�`G����P�k�[O�$@à�2�;  �#}-l��#y��X�׌rWȹ��>�=���7���%S���B��a�C���?�k�-��o �lWfI�z_��f�t���V�b϶Cn'�&0,�L�<}�8��84�]�������䃏��;jg3��5%5���ɤ�ʊ�?��ƴϧQ�,�����$�ߋ�2��u�0ESUW5VŞ{J0;~%�̝��i7��9����J	�,�z�J�l�
�wx��a��1�=ębt�t'`���p�귒J��_�yU7����R� M�v�I�����ao��u�sQ�S���;Gr�e�NΛF1X�{�Y�."�x�]z9��xo����l.�~H:%-�<��gR�G����'��	�F
���C�&U�,���U���@TD�1Jf��:�q�*��jFb5�}5#�h�z��y�e���ƍ�����"�������wG���T��>wt���<éG�k��?p�HMfU0���R�h�������+$�emu��1E*��:2��|+�Bq*�L r{,�G��
Z��ކ�(��k'���^�P��ȴ��01ʜco����<�.�1�q�˻9b+~HC`_��UO'���D�%8aCTP�x�V�&�a'�/$@����O�}������&r.��9vID�H���$���!��Tj/�Fٯ"�D��A�P��갞�mq�ִ:-H3��ϑ\���3]r?��_���9K����G.�v�H�vsJ�z�ck�9(;Pi�N�y��p��(ߡG#�O�v��0~��菏B���'�̌((��he$�-�Co:�S���	
 3�Π����b���<(B��_��b��tˇE���G���hUt��{�5�_������V� �������Bw҅��G5>E�A��w��W3�$����,[UN��qW�q�h>��7;iq� �6�3�q%��}��∋ڞJl������I�n�ę�����(�nY$9���/��V$�;�E9*�q��uX޷��a.���{}��:�^)~C�#�V����4Й������{ ~��S�q ,���l.�3c������{��f���U�����&�m�g�yd/)�'cH�I}iA6l��f�.��U����}[	S���$�l�6ߵ����i	0^/��{j�n��r��U����s�����aHDZ���P��)~���(�r����R�����Q�[��%� =���%M��N�_��y�Ѓe�����3?��!w�S�|p\?#����py-��\�)	@�;R?�LZ�8�Х6o���%8ؕ�%'�L����U�^���$6��(��m�c����sO,U��_�Z!ou���
�M��.U9�������
��Ǹ�iJ��«��vR"9@ȭ��T�����ި��R�.���s�15E�
�v��`����Z#AAZ�c��8�,�`霻o�����S��2g2j��P��.�(lC�M?�������M�5U�f�����6��=��q:1���h�=O�BA�$�&ƣ�[{���Y]��l6�|S�oU'=C�뽑k=���n~Y¾�#)v2�R��`�P�!�X|�"x�u���;q���*Y��Z�0�c�A���=�̥��ۢ��������ٴ&�EW�O??|���l�Q�B*AT�(�г¯d��@J3:�a�8W��T� �	m�Ȭ�HdD�!�P/������Z(�`�&�[Q�u��>�s�����S��Z���	�wϷ�r;&���D�l���?���i�L�8U`��_8,]�i#���r�yWr��6t~�\Л�-
�I���,eʢ�"��҂=��S/(h�J���3U��s"thI�����n~�G�uliЛv�:m�O��/E�M���eH|���d\�_��oF]�Ω	���f�����x4�UB��Rk�Q��	���K�����֛�!�2�a�;��C�ޫN�8R��P��2����#ϙ�Z��y�]�+�!Vs�T��u.�i�NՓ�j��K��s]�ͺih�'e��e�S̠o0���p,�	9�����P�{�v�V�KU�^�3��SGGB�;���@
h�S�v�Rz�cvx�Oyl�9��1���.�-p3 RT7Ғ��i��Y./�^��f�mkV������P��L���e��3;�wì�w�;�گ��⳽"�q��Czԁ���u�����%�=�_���{<M���g#s���E��C~�#�����N1��C7Ð�������@s�u �9���ٮ^$bQ��dlGAu���MM����_�}3��J�9�7Kn�9_'�ޏWV��� K�SL�" �ڃ"��ΐ���?� 

�앟�@J�y��9�Jj�@X�-�X�>`T��kd�'f�es����4p��uOi�y2��;캨����ߺ���Z#o�|��ߴ�ۅs&̇�]aŮ#��^P!8�,��$��1I�w��Qf�~�'�%��ϱM	����I�tl��e��_����0�MS��pqo���oi|��/��Т��V2 L�Z�G�̇~���6T��'�θ������V^�X�y�N�ܹxSr���le� )��Z�g�2=3@���;�	�,�� �����҆.>�>���įu�L.�ģ�%V�b���=8�(+����#U#�|�eٚĮ�yK3xOՁ����mi�5��uEu_>A��T�S�-��=��ˣ��jX�F�Dၭ�%h�������`��R����`�J1HO��8��JAˎ]I�	{Dg�����ůE{�MA�.v+㮈�W��� ���Gz�P�A"���6�En���v֕�_�j��U+|��H,lzO���-k.����[����*��3�����'��ޘ�T
���S���2���7}�j֋��[�$j�dO�֧�"e	������!���6��(o�:�]m�0q��Pb��%�k �@��=�mt��
~'�Ջ�^n�|�[�G����H��Fx>�E�%/V�������E�Q�6E�$���	-}�i
�E	�?�<�o�P����( E�c<��=��ڗj�i&^���îg�KF쇒��6B5��s�i�j>c1�� ]$Ԋ{:S"�U
��A'�f���*{%J�X�Řr3�`"8����A��n�sF���i)ˤ,���/�\����Jh9�p��ł��{��b�}�_<�'BٴO��򝁮R��istd�
����k���ԫc�G�-{�~'�ژ�ġ� ����.1/s�7����]�ơ.��jKz����/�m��@�o��yn��{���^^hW����lP.�.}��=�{��{����B&O�\x��ؾw��L�F�l��|>�LeIqQ�r�3��~�_ 菃l��,�B�x$:�E��?���-��t�o�j �fl�ϑ�DH����}��ӝ��y$�nR�P_���9�O�I��p�I�5#��Ķ�v����[Dea!��5 �]{�&l�P5<�B��p��osc"��K�����\�xChrфU��M�(y��ШUu�qYU9/����0a$Q�S�m'	�J��n"��p��~�eܪ�yn�1�y 
�𯹑�����+<	~:kg�r�
�B�Z��F��3��m�H�o�Ͷ*��XQ�7��3�$���Gt ��7G��|�7��6Q�yJ"K��ٰ8��*�];/���C�ⰹ:��Pxlʭ�'k��g8�sj��8��Vx�6a��#f2��!�����+��8�Tk+E����Ű��*�	�
,��0� l#V�q)Em�u�Ϫw���S�z�a�j�RD}�B2��:�m��j'�
�E�;%7�,5�H��(6��R�G9���/�����	̆,�÷����fl}�{.ǋF�^����ˉ�jٺ�!f������L�F���w0�k��?��Q{1/-#��HG���*�]�dm.P�-m5��8:_£eG�.�#��زv y�������FR	��׃�������=-14�*P��Y�V�2��c�=f�� �qW �u��L��(��"��	Mp!Iȫ�ن���vh:Q}��d�Z����A6�ڨ�c��M�E�"`��{�y3�R�Af��� ��Uƺ���Yyz�Б/���OIMh�w��������N%Y_�B�����ܼ6M���T�pXX{.X{t�b�r�N|������P�0�-c�C���i�����Q��gX�<1C'�d7v��l���tx�J���M�����m���l9\mp�����+2�]@t]�e��T9��6JaYt�;o*ՙ���>����$*ٔm[�+����
Gǀ���sYP�#g\+F�.�Q��/��F�ݻ�(�[�:��Np�I z# �s��^�<Q=}�#��ޕ�`�驷s��fRd���~�� Z�% ���1�ʲ��MX2Er�N���ޡ��~���B1�عЯ��:�I�k�8��<�P���h��N���*ޑQ�rt�J��y���;x�O�ϔ[s���6�s�@�ΝU�Q���~M_�^��mKk4�1Y��sE��K�@�hl��������/��Pz��3��Q���Gׯ=��u�H�>��"�h6E�5������V�8Xu��)��k���R�U�(��]O;���|O�����?F$>Mo<��o{�n�W�4��B������S޵_�n ��4Z8^��Y�f�ó�za��!k]���QE
:�L�Gl���\�B�~�@��`%қ�+&�3�V��3KZ����s�Ti��اK�����+y�3<׸~�Zݠ��B\A�>[�W\�2��X�k��\�K�k#ɑЈc�b�*l�B�D`�Z\�1�ʶ|]�4�L�\�Ɇi�/|$j�Z�������&Q��ʇ��BW��<���ྙ�Rv��te��6r�\�w�\���pއ��)oYt8<A
Z��Ѿ�ʣA#]�|�;`�󩨽�H^yBDC4m����yL���5k?��h+�u|��x����*ػ���6UY|~�SVf�|[�&��Jz��T�`[!�}�Z"�Bn.���M��9�/w���i'.n�Mt�PB$p�NG�kي;�@��<}�Eh�S��@������( ����C~�Y-;��b�s/ΥeE�,��&o�c4Z:-Ƞ�*[�H|�ſ��%�]��S�)��D:'@�,�gg�xxZ�i|% T��n�@]-[�ܦهA ��K��K�4�<C��gK��?�S3����|$Ӿ�0Md�'Z��`�����V�c�e� uZp��P�/�@M��>o�d�=R��Ƒx�녈��*��`h��Z�&�w���:԰�R��R�_p[	�>��?�gI�������(RG![]F�:g��H����6��do3�q��J�|+=�L�������dW�����/.*|��Zִ^��7��.,���N8ģ�!���u���B��w�l��L�
2���!C�7�J��cTZ|���ف���J=��[AI��*C�d�?��T���A��,�̩Il��ig4{nו�r��Fe/H��jk��<_�ub���#�T��~���s�ˏa}V�0�Al`�l�9���C�3���g��gr'��r��1�j��\/H� �\���T����-�Z�<�v��P��W�j�\���?��
�
9�oRpqG�T�7��q���>��:%�#@uȈ�L���a�,�,��}��r��R����׶)�>�4j҃oԱ&¯#�xl����J�����;���Li+
S��w,O�P4:��x4o���M���m��/2zɕ_NHo|���*\���S��\r~�,�C��D�0,��d�Ci�sKё_-L#�_Z��Syp�i;�] r�L��è9���P[&{|�Ǖ�����՝	� �����u��KNA,����EHwwF��
c	B.�
�L���>��`�vO��6T�,��ҳ��+�%�9ɰ8P/ͻ�ʲ@�;�
�9��gq�����fF�B���+Y-�烉Q�.��[���6��׎�l�n?_ř���9��el���}�bcSӪ#�I*�)�pr�k@~oO��B�<B��m�a��Y3?[��5º%���*��%��ss�#�?��@����۾�['P��}�V�vr_l�	َ�3)�J?�3hP�Uat	�h쾍��Vc�R���*�MP�AA����ԯ���G�U������M�8�7}��}�'�+._�Nn�/s<��L��O!}����<����2��������ZE���� :Ib�� ��9�}����<`�q����9VA2��疽%�n��� M
�r���w±�p���*�Z�q��k���kS`�6<����r.$�U�F��Y_�h����&\�+	�] 9v�

���:q�,������D"��o|b� S8� �~[��S����g;W��H'�=4x{|��-Ц]j�P�0�Aepz�B�+H�Q��t�&��wb���E���g��t��c���!}�qGJ�Lz�.G٫`�m-+�|%z����/���R1��j�/٤Σ��G�$6�0k57`��שm���O�_����ZX{1e{Y����R摢��[������q�e��e�YH�E�^@���k��O�����
˿C�%����9N��j���xv����mA���i�?l`�A�����ieJ{`w�Ӌ����f���j�X��6��/mx�V%}��`�Ƴfg�c���w7xĜ�[�����5��T3��"�g�U�,��/~�����p����m�'�����/z�׃�"?d�8�'OVR���\_5]A�2��4�b��ߛ#�+8�(K������m��lb��<��'tCGd΢��A�*���[�*�"��ܦ}wV�D� �a��c�619r�"��]2�� 	\�U�֬^R����z���������F74e����$m�O$U�����Ɇߊ8���Rj��\w+,:���1�)k̸6� !��O��%m��T�!?��[��im��?D��]���6�b�b�^��:}|��c�C:��}Х�aO�Y[m�k����<:Q��AZ��я�>�Nm;Xg�9�妫�	Q
���o�/ܺ3���Y��G��Ѹ`��ߊ��������!xo�qe�lt����9+y���̜_�4S�%�v(��������E��`��Sꚣ[�j|��F�2Z��&
��V�S+��� ,���\�rK �Q_%2lSCv��2�SL@�������m✾�N��
,�&6�� �X�_����w�Q.&﬍�{�������Xh�(m>�@7�=�O�.��J�IX,��ő��V�^�+N����Fl����~(7����u��Ov�_��$�*�a)�����Kd�,�/0�Q��Sa'ZLCgƠJ4�q%(���lL-p8
R�|�7�H��^1�V���[o��O���J�~,Z���a��f��sA%ƴ�%��^+��\��f��U��I�E��-�HTTt����\qQ�X����5I��l�7ε���b�Axu�
����A�a���\άhVifW�u �K�?W���ɧd����Ra�
��lg8Q����I�!��r}tdG�@
���9tv|k�:֘��{٬s-7�͋pv�U"�8�54��Q �Z��=�\.�I��܇�p�]2�sЮ.�r3(w'���ǟ�-�,)6����IN��{w�K���ր"��Y�8�n^�,��˕���MA�����'�q������Nr�,Kt���.�Քݣ꫟\�n�&����n�h
���3��� }3S�����Jɒ����Tf�B����=�w�L��Fρ�¤c���Dzݴܔ#&F�h���ɜ�D1��K/1*�0�d���`��?�rA�b�)-jy��?4���>�JX����|��Sw$q���������I�FO��If�t������{�#���9�/����f�k���ѿ˸<�Ih#�.�݊��%��
<�i��w��I�G@����ڜKƣY�ܕ�O��}C[Ţ��x��d�ޓ�5�=����k�6g]�1�|;,� �yak�-2�o`{@դu�x��]~�o���gLe1^;ex��LƗ̺TsQ�˹ࡈ�MuY-�Sz�"'�ǭ��
+�a|����Vl��)�V�.�/�!�^`L�7.U�wa쁅O�+����}����G.	3�pn:�&0��ѐ��Qf��CG&�D�\�S_������Uf�"�1M-c�>"��q��A�Qp�mOA�V�%:8!#O�ށ�"aa��)��Z�j�Bt���G«A�c��i��db@I`����@7rLuʘ K�f��4(�* T+�r ��d]h����lE/����Gֆ8*8��Z�[�+��@�}s��~W�L���O�9Յ!�){K�*�O��ˮ3��ji�9xM�ei�ؓ�&;ہ��i��eb0K����V�ڰ�t�Y�B����e��j���S�����:���l�b����P���Θ��`�F���7�b��&1K��-(x��	�b+<-�$�Od@j�w�G;�,���03��	�*֜fQ��Bw"(�S�jb�$܈pR��7��-.b�iA��@=ka��8���儠0���֐?�2{����~d����FJm0~�͑K0�߀x�;�*�ߢd��<��d�/*�C�ű�>#٪�=�Je�w�6]��j�f�I"�e�
~�6g2���e_�?�Q������N8s,:��C�����ol���c����O>!a�s��!�0%X��3��r�a�.qhǺ>�Z�ҟ�`��	� �TG�/����2X!����8�%/�]�OvZ��Vˣ�����YAg�F���l�v���vfv�.a`��@O�|�ODRs�������V7]���⅓���Ш��q����F�=?	R[���?�ĝ�Ku1��w��?�[�0�� .�