��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR���b�z�>}�����.�z,yN<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR���b�z�>}�����.�z,yN<��;��� B]�pE���	x]̃Dj#^Da����M�Ov��12È�pT�7y��z����)�,�˛D��w���旴4�����:��@���b���$[��-�4(_� .�4TM���.�a��jǎX������n�q,��m����Zߧl4���0�?�1~�x�cq����Us%�ꤸ�����%U��0�$$� d/cD�#��x�۶�kv�+3ǆ/����`����ǆ�$�"lj-*�NB�悑/�ߘ��~�eAc��o���0��H��k^�;��;&0��\ D����M���ѵ�Th�fܯ�ko��^]�����S�~����p,+$\�M�T�d�$�u�}�<��O��<$e|����w'��1�:�Ω�[@�qR���b�z�>}�����.�z,yN<��;���u��w)�S �J���vy��e��m*q;�K?���p��O��Of�+���jv���z-&)�SD�:�Ä�����N�v����
��e��o����1�����(��^	�܍�1s��i.o�*nŐ�u�l��êME���W͉A�?����i��vp�$_<n�ȳ؜k`��Z��L�R�.�$m>�-�_]�og�]�n������fxQ��)��\�4�s�gD�bOq������ǃ�8ƶf�,w9������ֹY���8C�j:`d!��tW��] ��[+�c�5���AQ� ��_�^�r]��K�X��K�zb$z{
� �AH��T���x�3�Z�<uo��0]��;�*tD�>;�L����� ���>	I�멲ٰ�Ř�h^������*����	~+�<���p2��O�_Kc�[_H|�eĕo��tW��] ����&�[>�y��W�y��MqZb�L� �k�#�l�w|ü��}T��X����::R�nҎ� ��k��_֦�j0V5����
� �AH�h	_�fx���Z�<uoz�!Կn��i}3�L����¸
uy�BU��f%%eo���sp%S�y,Y/�7{'3'�`�m�!=�y����h�}K?c�*�S�\�l#�+ohCoǬ��oB;sѱE�?�m��l�j���N�=�����q*\�9X�����XQDi����N�v��<���P���d1���P��)2R��DU�AP�nJ���_U�t:�W�g����J%�hu}�fO`�|�2z�R��톋%$ n��c_�Jh�5L��p
� �AH�+�6�O�_M��RwM�麶V$�(k��n�L�����r���(�����5ʦ�&�d�I�_ K.u0�p���?�o�3�P2G�e��-�u��w)�SU��T�d�I�� ���I�"{��&U6g���Kf�+����Z��r��p��>����}�F��qt4$p�)�����W{��!�*��x�6p.��k�8���҆�|n��tCP��뚽���I;������4I�0��U�)�(27�׳������<�6�+r
�M95��v�7����}ʬd�ŷ|�v������s��"q�Aj��6�T-t���S�X��Z�Ʒa�o�u�/�|?F���DB�T���xĄ}R���~�$�Z��ДJ��_��"SӠ�|&�:h��_���&Y��V�F��2��+��T����5yi���FnBƕH�N�4�T�f��Wj�����gB����/��PJ���9� c��(�U����	x]�W��r�B#��ئ^��B��gF�������8e�S�O1���kz#s*�[A2B���d9@:��'m_XK�B}��%%��T�1
��Q���+�7x�Ym-46���RL�a)k=�c`SWH�~篟|�>�w(�ոK��4�L�9����E�E����}�c��_�+-�S�A���T�*�QKUY�}�h<r�O��C��0���C�f.�j��r������5�ݍL
�tu�OMp�0V��]��b�4V�U��}~d��w-�c��X�X�;��@�b�A{$��ش�Խ�ã�E�+�iP[4!{���V
�:/YD���RL�a)\:���}��~篟|�:�A+�4ik�eȺCs9����E��j}g��*�>�i�$A�8'�+���w=�:<~گ#(n@��\�4�sP&�O�S��Z�o/5�������y����E�ЌֹY���8�'�-��p�~�@#�9��Ѳ>�љ���>��+�q�������c� S,?[
� �AH���<T�%4M��RwM��#�r�N�y���V͙�L������ �x�"ţX`��_/Խ�ã��/5���sӌ���(�u��w)�S��X3�����:Vx�p*�Hؕ�(�&㪡g�f�+���.I���C=E�o-
���x��-�/�ˌ��D.�1�M�w���I�u��� c��(�U����	x]̫f�.(`����7��=Ru���p`��S�O1�༨`��*��½<�!r�O��C��0���XϹ)���J��e4oDIA��{�S���D	Ey�"o
��qt4$p����)�j|`�� �V;Z��&/`�r��Z�r�r�Hi`'���\�4�s�%�{�[�K+8�M%��s� �޹ș���ֹY���8
��D9v���o}B�,r�O��C��0���1��ǉ��s��M�F��I��k�i�DE�AjA��j6Y�T �����y;�j��-=����Gq/x����n!�z�BV� ���Y��ƴ���(��}���W��4��n�b��k�8���҆�|n���.�hg1��fY�?���c�t���U�)��:���[^=K�03�>	o��\~K�f�h�9LC=�`���l�����~x�k�/�x�˳�����zt���:g���8�_�uf�����;t>
r�O��C��0��#}������d�0�j�h��p�)l���AEP��]���_��݌Aջ��b�țQd���O�O�����q��hw�s�͹m�!=�y����h�}��[䁻�(�Y���mE�ti퐴���B��0L����¢��~g�Dm��Pf�
� �AH��KH���(�Y���m��'��*tD�>;�L�����U<˝�3%�
�� ��`C�4ː��c!��`�u�Tg�m�!=�y����h�}�G���Aj��͹!jr�SAoB;sѱE�(N�ᜨX��eʣ͜���_tKr���"c]IۯWW)��j)yc�n�.�_�t��|�$J�.sF.g	܉P.!܃��L~΄gO�3'6c�f��7�F�����,6��Ū;`�-�[[�������y��hH�r�Yc>U~�Ƙ3�q��k�8���҆�|n��1���N�Ee�Wj�O(z���x_��U�)�w�����z�\"k]δJ�����?�Z�cU}a�F��R�}vJ^fN��ݶO�ذ2�����;%��7&�r�&U������G|M��W�J�.�m�!=�y����h�}Jpv��ư /�1�Z���m{�>��U�)��+������hQ4`�����-�\��$�Ff��u��
��u��e���ȭ�w�^.��]�!{gZ�f5w��jJ���_�wl�9��v�����1���
!�~~N��	�Ȓ��O���(�Z7�}�!�k�좏1Y�� g��N���RL�a))�kc�߇�K+8�MIWa���؉$|��x$ֹY���8�
��c����������z�L�2��~jV�F�zykR�At�r�O��C��0��D�[T�Q~P�O�#��V�x�FoB;sѱE�q��_�}eO��	N)�`Ñ�ԆD^�E�)��f�ɨVu��7���	x]�fX�eϝ(���� �h�ǜܖ�u8t��Y�*�y{�NѐR"~�u��w)�S�3k:�(�-�~篟|����T�	ءc]"t�39����E�k8�Jlk�#�(�\��wŷ�8�2o��RL�a)ѻtUWR��K+8�M�Mf^HB�Lt3�T��%ֹY���8����7�R^�����K��',h�m�m�!=�y����h�}ILhqi�{�k6�����c��C��3���U�)��#>fS�H���zϻ��2�v�;sۀ7���\�d���|�;ܡy�`N�z�������# H��9%J��!�:e��x�,`��O��2$6�sI�A|����T���|��W`��>d���WM�P[�������*l�
� �AH�}��� ��>,�
w�?���w�F@Q����{S�O1��9@o���'}�._�+��m�!Z�TH��RL�a)=�y�~ ��K a[��2�O3�ߵ��N�g6��ֹY���8�SU�/�.JLf�d��"Aw������c������bj���2�}�����]ظY�� ���A�=��L�̙�J����6�m���Y�8{�|�a�.��"�U�����;�Ӏ�p!!v*!���e�A��r����$l��ȍ��б�O�F�uw{j�$?�ď,c0�2��wv�<֖�����E�q��P����t���۰D��"�Y�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��He����L#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U�~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�ĲW��,)B�|aڧ������'SR����.�}|��ι%9T��7���S5H�j.F�YZY0@ìO�tw:g+��T��٤�2[51g.� -��E�I�?g�f�$��P�`
5��*�z��Yk"1/���qH��^��+o��	g�y�+��T��٤�2[51g���i��T!ea�8���*���g S�ĲW��,)i/-�#�~09h�i�k1i�f1?�e�Bw�M�?_W�\I���A#|��[�m���w��L�����'�@���,������0�ea�8�����B}rs���{Z85۰���N�l8������t�iZ]XF�@�ú�Q|��7�ǋK=��ͨ�s B�8,?CmYz(ݲm@��w?����+{ߗ� �#O�/�Qw-1�=�p��'$���Ԫ�3m������D�[�8L:i���İ�
��E�9Z��XON&~}�=Ll�����&}0�@����OYd-PJ���9٤��H�&�&l������ nU�IÙ=�Hz}��u�����\{F˯�+)���u*K6HT�����N�~ `�T�v��1���;ε��IÙ=�H<z,Ҽ&�jV�{+穴ʐx�?�'n�^0o)�X��2S-v��B��q�T��&�����-N���\�v��wc�}�![��P�ǍZ�J�����+�'T��N�ǁ�f�TJؓ���!��\�v��$DJ�<L	�>���Ww�k�̔`N�����n�j�Q�����d'�'n�^0o�!���!������"�=b��v�8:.��w���\�v�X�zgq�鄿0O���ġ��,��u*K6H�q	k���A��2�F�PY~�y�����[�JHn��z���G7�����o)�]rx�y�Zgl�.����JHn��z�Sp�}�f�HfCf�63���ш|m�Q� �٦��dk�r�&U���0��PW��u*K6HT�����N�͹ ��I�Q4p�/Cj���C�1��;�׊�:zL͊�q���\��;�,��yN4&�iq�VD�Lg�q��Dv;gJHn��z��r9�3��lT7Y�PG��l��3\_ q1j�iϽ��j�Q%��{S'��{,�
w��|ݔ�3�5�}�]���x�]�V�����Ү���/^�yQA�?��{m����
q<O�A'�u���.���hGD@�F��q&�G"f�x��r�Ti��7݊<Fi"I��ao.\C�k�ף�D�~4#C(�}�IÙ=�H4��%�Q��B�"}�fÁ��/��F��H��\�v�[�w����)t�O9�1.A�3q.��
�W}L���7�H)C� `A��~E�.���hGD@�F��q���i�����Y�V&��A��.D�.���hGD@�F��q���i�����Y�V�~G������"�4];ˍH�cPm���,%��\D����ά�.a�*\�9X���fˉ���Q�Q�q�o'�4];ˍH����������bJ���I<��fҾ��9��ЂDa��(o��0��7��|g�Y�'���Xw�f�VHF��Q�#<4^�v�ј�"��Z鎬����F�71�B�������%�N�By3��<�]�!����M[��Ǣ�L ʞ��0��m��x���j���0z�cUL3�X�j��7$2Ӕ�1���_�wa(􆿳�tP"7��%e��0�U+�qbp@��wbk�$���7Z���(�
t�ژq���U� бb*	��|	�WI�����
L'���Xw�4��}�<�=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ��B�m��U�;�j����Y%T��BPe.��xu	�L$�����/���iP1i�Q4�x#�+�B�&�g_�
�����Yl���#�]�!��	Ǹ�y85��(�C)&���lC��U�T�\ �͹g}|�H���p��b��e������]�!��	Ǹ�y85���ǳ@�M�H�ɇM��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+�ڔ�wV���C�Sy6ג��̹��/R F���9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8�����B}rs���{Z85۰���N�l8������T���u�I�	nrB��ZaԘ�������յ�}$|~ïSup�xg쬉� }���n4s1��7�癆cg�!������:"�9ʮU:���s:��t�5i^��EQ73)yn�w�x'���Ě���aT��3G��?�#M'���"��y��6��S3�ߟ{����c�,�V(��_�8)$���}6<6zY~G��A( ����_ $}��}5Xx�	�+�&I(&�L�ӵ��)���>�ѻ�5����g����ĳ��2S����"ܲ�����^Lma��C�<�Sm��q��Gh�3�!1�F$f��_Ub���uQL+����6��S3�ߟ{����h~E��+m���L����Ҙ$7o4 l�5Y�0`�WC����B{�LϬM��+��!WS���
9Wp��� gؓ��')-W`������a�"�fE~�cb�i0[����8|��`��W�U	EX͇�jO���a��Ó=�vzFg>"�vA��K1P��)�b���g��� ��"�~�>����;�P�t�5qM�4��o�Lѯ����Qٯ�b���L����Ҙ$7U2�h=c�ugÕ�KF:����Į��KH ����p4c�.�U	aw����Ѹ��ln�~8!��vp�o�6��aH7luP7���8-|�DF
�j��6������1�R+-h]�0�tW	�pg^��Pv�
�\� �jO���a��E�' �!��"� +}Z�"��%o�&��cay�[}�	76�&�� Ӗ�t�t��"^��#��Q���@��q�r����開s��m�z����9C��,ў1�ˏ�~ǹ�z��hbvk~�#x���EE��n��V����#���F�O��$�}$|~�﫞��fS�Q�S�T�=k�Rm��̍$�D�u&g()��ikp���H����-��԰�3�#���F<�X��j������&<v�}����1`�O�t_)x�?{��J�SqVEG��5���-�;���N��}�!`�������a�"�2�ʏ�"�<��E��b���a.Y�wg������F��O�z��K	pgu�5T��$ VRMR��,�*�K0Wi�l�U����;�� ��-�3��&Oa9Y֪{���ɖ?��_T���a�aq��ڷF����/woP}[�.ᬵy��5_
� �����3���ne
���HK�0,���U<� N��r*�jB�B[�)x�?{��J�SqVE
7�Ԗ�E�.ᬵy��5�H����;���<@�� Suiӑ�xGe�;���N��}�!`�������a�"�2�ʏ�"�<��E��b���a.Y�wg������F��O�z��K	p����)Pg�ŉ�u��M�B��{���"���@
H$��j�>���?���B��Ul�~ǹ�z��hbvk~�#x���EE��n��V����#���F�O��$�}$|~ïSup�xg쬉� }�=k�Rm���ӑ�xGe�;���N��}�!`���Nj�a=�t[a_�?��J*�Rs�0c�툼��#���F��3�k�n�V*ڎ�0���J�և3
�v�v-}�	mp=b�ɝ:�3GV���J�1���-�".Q����>���?���B��Ul9��f;���"��y2�LpOJEl��Q�P�]zm?9ۄ��d1$�Q�<om���b9���M��A���va�{����U ��z�!e���im�th�U�CLB�D5�O�X��WG ���y�9�3��4��A�(bGuj}��8�,ԱvD3n�x(�i��/Rz��K	p��ay�Ȇ^���x�k]m���C�MV���%��b����3X����a�x��M�ݭ�~r}*И��&�������Ŏ{�"��}�偢��%�<ͯ�G��R'),��`�@ux�[����3���ne66�v��G���V>�R< N��r*��حFہ֥��ع��8�b�R$�Տ���i���a<�*^e��J�v�t��Ʊ�_�eD�I��3��oE���$�8@�ɮ��U���#Â��&?��Nj�a=�x^1⩠�^!�<8qx(�i��/Rj���;��D3X����a�x��M�ݭ�~r}�֫��XA��Gm�o�j��`KL[�{W�g���F�i;�:U�v�3b��{"���,���"��y�xI�2^)b��@ŋ��5k.'C���Y�V������p�0ty�P���Պ�`^��3�J��\�v�w�?�b�>޼�\�vř9���=��\���.@A�-�]s�(_�<�� ��b�FP&����҅JHn��z���������x�&�F�]:��='����R��e%�2�ͼ���y�]�F�D�+�:�G�9�E᭗��_��&Yd&�j}!��n�͑��LK.I�:���3k��g1�e%�2����莇����_����~���i�x˗9��6�8�d^�ϓ��ͬz�Ť��xI�2^)b��@ŋ��5_@&:������;�R�I͗� �-�`)��\^�#�f�R�I0���ԏc�r�(���JHn��z��|/��N��hk��Y��A�m�(�b9�����閝eu�m&� JHn��z�w�<¯�����v�8:®xԜ��H1Y�ΊS&h�5,Wl�/�O'�=�ƣD��8!��vp�P}��O��^��mi9Ů���z�jaV�,�&{�zYa䃾���Kl0��F��j!-`���w�|ò���
��_��������[a�[�J���6�@3uå��:(�
�*S�#���F)�S������4���XP��ȭb��v݋N������5R܅dJ�A���ۖT��Go1z�Ů���z������e���ݟ���O�͛PA,qLn��S�W�
����uK�r�&U������G|M��M�~}�]�+U�HJ�h<��}@�ͫ���r�3�����!%Ah�%4
>�(_�<�� ��b�FP&��獶���_�(�X�)�v�V�.��b9���.M�"��Ӗ��s��2b���!h�b�TG|�w57�S��pN��B�)Y�+U�HJ�hn�./�������|I1=��%Ah�%4
>�(_�<�� ��b�FP&F�W�1'����
3��FZ�ޑǇ_���˱���v�0���f70���!�`�(i3�����5	��M�-��#�g#���I}��NV�MO���9�<�!8	�I]��� N��r*�$��ûX��kRCլ�����`��&f��w�'�?t�kJ �&{�zYa���<��ɢ�U8��ّ�k���H��@!�#-�[ҭ�g���y��b��v݋N��������c��>z�Vg.N�������6���|��"5�o٥۪	�}a�iQ��ׇJ�	�LÆ��/�i�����܍w�S}9g	���W���b���p��=�^���3
�v�v-}�	mp�����2x�N?Dd�-$#�0$�.�-v�Μ(4���Yk˃Tc�δ�0���'?Rg�\�G���nQ�rV���1���X��WG ��D����jF��b�(� �	T�����3
�v�v-}�	mp�cA�N�Y�74��LM�(�� 	l��lBýO����ezꥦ��r���:�����C��괽���5%�"|R��9%2�8���x�Y�1G�Sזi�)x�?{����ҳ�ET��o*|�[3�^�P�qjhbvk~�#xe�����t���3��Μ(4��fU��S��ɻ�7��M����v�l5��� rư1�l�_�4��׏�����M\]YD�^�O�<om��Ts��E=�!�Wƞ$�FA��mӡ���<K�yw���-�3
�v�v-}�	mp�^5��$�9_��i�D�,����3�<�:@�@��\l�垹Y8��#�8���w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�w��AW�Z�y��l�Ow0H��G��9%2�8�Κ���@>��nQ�rV�����J [ܰ1��?�shbvk~�#x=�;����b��v݋N�������0'n�ڹ� ��yo�}�Y�PX�)��s����A���cZx�.��8wCc ,P��#��\��v�8:��MWU�?
�5ߧE4����{�A��3D�� <(rK�� ����ޙ���9%2�8�μq�T�<������t����==�x�Y�����5O�r�����Tb΃l�����}0x�PI��e��&�'��;���N��6H*��l�A���ۖ!���6�,N|��|(F9%2�8�Α��H����ָ������%N�ݚ������	5sJ�J�	�LÆ��W��C�܍w�S}&��|�7���Ɵ$v}�S滑���f�� ����p��}��aq���g0����Xjۙ�)��s���#Â��&?���J��6>�2�q�]��x`��:�x(�i��/R1`�O�t_)x�?{��J�SqVE�e�H:�I0���ԏ����[���Bf��0���f������C;�,]�eT�n
V~$�H�*x����=��:�H�*x��1d�ެپP۪	�}a�l0� �A(�i�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��n
V~$�Y���� ��@s'R�r���t;\`�r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�ܿE�qqRmF܂d�ۤ�m�>!��bT�$&�fe�X����)ͶG�q�5�
p��r%̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-���Y���� ��@s'R�r���t;\`�r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�ܿE�qqRmF܂d�ۤ�m�>!�����4c��X����)ͶG�q�5�=��ﯭk̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-���Y���� ��@s'R��E=���r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^��o�������|I~�I����uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#L�tD:��@F�W�1'����
3��~�/:���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��'#���n�{�X����)ͶG�q�5�	`�/��í��H��@!�#-�[ҭ�nɦ4��De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�O�β\�{!ˎ]":V���"^Be��Dc]�`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B�鉞(Q��;��b�=��?njS��}�vo;��|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*��'�/7Ii�^�Ax񣘂D-\`��EW+GE�Kf
�f�3
�v�v-}�	mp˜�ķ_�L�b��v݋N�����6�pnWwщ�(Q��;��b�=�`��N�G�g�r �����=}'t<��ġ��,.R��д=|��(Q��;��b�=���N��/*�A���ۖ�ꉴ�dyi#nĖ�*i�^�Ax񣘂D-\`�����SVc�Kf
�f�3
�v�v-}�	mp˜�ķ_�L�b��v݋N�����6�pnWwщ�(Q��;��b�=�
22x`8y8�g�r �����=}'t<��ġ��,.R��д=|��(Q��;��b�=澖f���e��A���ۖC=4�a,�n
V~$�Y���� ��@s'R�r���t;\`B�R���>_���!&�+��h�G6SX��Xjۙ�)��s���'��m�xl��(Q��;��b�=�ύ<Z=�	��U=��G>EK�� ��Ut�\��Y���� ��@s'R�t��&� ��"L?���J4[���w�����1��r�.Gb�TG|�w�q-2�;�"�2�q�]��7�H5�RF܂d�ۤ�|��F��ڊͣ�:Y��Y�^�f�s�tG�ه� �4�<��U=��G>EK�� ��Ut�\��D$��:��
3�t%9��&����1�%d6c�d	�Ȟ���p�o�QM�W?#<b��>
rw�&�z<aSm�6��`4�04�jfh�x#�L_����	�r��9��o���>6�P��%,��7n������A�9�-���Y�f,�s��Zrt�\0�{�q֣���óM�˄NKYi����L;ø\����?v���=!ߎ�΂l��=5;�D|�[�R�n��V���|ò���
��_�����,fF�7�1Y�ΊS&���0i���7����NT�<�*�!g()��ikp���H����b9���ʵ\���Ex�y�Zgl�[��j/Ҥd�X�VM�����a�"�'n�^0o.�ؙ�b�Ӧ��9���I5�4`UV#-�[ҭ���~����'n�^0o��N:�@?u�hk��Y��A�m�(xE8�ELE��&ċ�;���.{2Y��{�3�P���ġ��,�Q7I�2)��\�v�#�1�N�_�n�To�[��8-��-�3
�v�v-}�	mp��T�����,�v����f������C;��S���'n�^0o4��t-s�e�J�Pn\�H�4I�B�������y�r��VYW\�o���*ٝ�/�K^b�;��	+����4���XP���3Zk�E��% ��q ���h�c�M���v�8:mvvb��_�.ᬵy���=t/��g#������a2����b�������<X�l0��F��j�?��;
V�;���EWrN|��|(F9%2�8�������JHn��z��o�RO�v0I��'��_�(�X�w���vc�f70���JHn��z�9�Wz��
)x�?{����ҳ�ET��o*|�[3�^�P�qjhbvk~�#xe�����t���3��Μ(4��fU��S��ɻ�7��M����v�l5��� rư1o8�<����;���EWr��$�J݃����t����FZ�ޑǇ_����'W�=�-��/�D�ؒ��"��KH����t��(�z�=�j��\�v�Џ�I��$��cn��>��u��j�E��*�j�H��b�(� xܟ�,3JWA�%��fOX�����̏we ��g������%ng ���3�ҺIÙ=�HM�f�<�O���L��^�
h�tG�b��v݋N��������2����hk��Y��A�m�(�{`x��%5[��	=g()��ikp���H����zY�l��R�}vJ^��l�|- ��b�FP&�q���3B��*w�o9@g^�J<�b9���.M�"��ӖEKM�yW�T�s Wd2U����v�
����4��(_�<�� ��b�FP&f�%A�)!�`�(i3!�`�(i3�b9���.M�"��Ӗ����������
�x�w�������������� �1x�itLd�r:ha3B��*w�C&�5,���a	!33֬�lPCrM�Zc��~�/:��ǆQV���Ҥ�������|I�W����x�A/�n6�r\�H��/Sg4�y�)@��]��0�ȍ�x�>c�K����&&\�0���eYk�	�yOx(�i��/R�Ȟ3I	��.ᬵy��H *4�ڮ���Bư��9%2�8���x�Y�+���]���J*�Rs�0u����x/��'�ĮpYÕLM�(�� 	l��lB���U%�p�zꥦ���i͑��Ԣ���C��괽���5��g����;���N��-Lk���ޟy�K����t����==�x�Yu�~����J*�Rs�0u����x/�'��ޙ4!ֱk���p�˳c��sCF��[ S��x�%�/�d�"�hm�^�6/
��VLM�ǩ��8���׷y�S}m� 2�k#ʘ4��\��sپ#�J��v�8:I�}-��^R��	�ݑg()��ikp���H���ʤ4���aHUv�׿e\V��/��x�%�B���vs.�^�6/
ڌ����S�|���#q��iQ��ׇJ�	�LÆ��/�i�����܍w�S}���d����_�(�X�<�q��Dp��3
�v�v-}�	mphpL��m�d������g()��ikp���H����-��԰�3�I))����A�m�(ą���P4�=KmS��3D�� <(rK�� ���$!��8f�� ��}���x�A���ۖ��P4�{!� ��3�F��Zr�Z��T۳�͕��w0H��G��9%2�8��!����&@��(+���<om��k%-uב8)x�?{��偗#���\ԍE��C��>CR`�y1��r�.Gb�TG|�wA�2)q��FA��mӡ���<K�I3����b���z�òr0y4{�H�a�\�#���Fq������n
V~$�H�*x����=��:nQ�rV�)�YBa�g()��ikp���H���x��3�Y�^��q,u;�B�R���>_�qЕak֕��A�\>W�/Z�������u�`��3+��f������C;k�k�)%|�	�Ȟ�����hLKWX��WG ���
�����w��r|��߇(���л���.Ȃb�����V�I�e!��nH�W���:0>��� Q��!$�2�q�]��wc�}�![B�R���>_�?Iߕ��1ҙt&H����y�]x(�i��/Rh�x#�L_�h�:��p�3
�v�v-}�	mpҭ���^���b��v݋N�����6�pnWw���z3�:��c��%2���ʏ!�܍w�S}&��|�7���Ɵ$v}ֱl�40ߏ3��#Y�r/��5Տ4�04�jfN��������KG�5�zU��آ99BI|�6|����J%�hu��y�c�i������b?�*����f�����"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�t�%�(^?�f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#�P9(�bC�3
�v�v-}�	mpҭ���^���b��v݋N��������;B����z3�:��c��%2���ʏ!&f��w�'Xv��@�E��`;�nQ�ǅ�a�
ȍ�F�]	
~ao.\C�k����|�i�^�Ax�6�װ���='Ӏ�d&��(Q��;��b�=�OcDb==�7��%��Gy�ˆn����N��+�?ݨ���#2y�Z���7�A�6x��iY�g��ѵ�"xC��-�T(u	M^)FU9����g,Z�fg�4���R��T��̪mMUt��!b�4=y�(ͻ� ���7���ìL��-)6�oȔ�T�͒�H��@!�#-�[ҭ��:�*�3������w2}�<��bd?�&���u�~A4z��4^i�u�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�q��uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#�g�r ������w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x������|O�\�+�q�� 6x�@TW1R�X�L�tD:��@|��������2���t�I�� "\�H��/Sghg�R~G�����A��%,��7n��̥��}20����9��F܂d�ۤ�����ms3M��o(ͻ� ���7���ì\��2l����Q�=ؗ���`;�nQ��A@��sZ��o���*ٝ�/�K^b�;��	+�/��~�;1֬�lPCrM�Zc��ʪ<4 �"j|�S�
���N�@E�V)�jP|B�1��6�G۽^�w�򪥃�n�{��l[hbvk~�#xM+)�C%�&|���BY��l��=5;�B�8��\]s������&{�zYa�k�f}�Ɔ������g����;���NC")t[p��]s������&{�zYa�f���%��)x�?{��
0#`�1��n
V~$|��������2���t9�'��_�K�z��d>Q���G&o6��~��<o��!h�b�TG|�w�q-2�;�"�2�q�]�>��O˻����|I�w�63xHl��7=�[G��"xC��-�T(u	M^��|A�IU���b���"~6���aq���7��Y^&��fx'v�ao.\C�k�4yn����q���3B��*w�������(�Ae�̃B���K�<om���м�1#���q���3B��*w� eY�NA�J*�Rs�0$�9͹)��X��WG ������*��P3�lWD�q�5�=ڭ��"xC��-�T(u	M^ �(팵���$�J݃����t����
0�@lJ*�Rs�0K=X���d��h�e��SV�Cagi�"��(Q��;��b�=�U3{����B|�S�
���N�@E�V)�jP|B�1	S�%̌��n|�
H&b_�n�To�[��g���a��>�8-�ށ���
3�E�ʫj�>��O˻����|I����ZqM����
��\�H��/Sg�zH^x���r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^܊@3+'�tL�a.l�n�)^��o�������|Iܲ��9m����͵De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N�����K����������\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|�zYק�̒�H��@!�#-�[ҭ��F6q,/̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t�h�N#�Ǐ��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
3�м�1#���q���3B��*w���k�t�f��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!r�
C���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g庌NA(fۉ���$,��F܂d�ۤ�m�>!����J�Cp�������s�`�|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*;̊���z�1[FQ������-K��s����M�;䌚"\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|���sHT�f��H��@!�#-�[ҭ��F6q,/��h�`N���V�I�e!��nH�W�l,ѳ��=c�f������C;��?��QX��WG ��BE�r����`;�nQ�ǡ2�!�7$��q�e<r�4^i�u�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�qV����Eˎ]":V�C���*DwS9<~�p_�X����)ͶG�q�5�SU*�<�)��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!v6�RMS���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g�n�J+s����$,��F܂d�ۤ�m�>!��˯����9Ǖ��A�\>W�/Z��B���[@���[��QPw��r|��߇(���м	I���������)��H�'J!0��A�6x����V�C���Ul�ٻܔ�ߎ�
1y�A_`OT q��Ko.g()��ikp���H����-��԰�3�I))����A�m�(�A��PmP	�Ȟ�����hLKWਠ9V�-^֬�lPCrM�Zc��qP�U�&�De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N������ᴶ;R���F^GQ!�сn����+�Y���� ��@s'R�Rw�)���$G����N�����,eS=�oA��$�J݃����t����9��b>��X����)ͶG�q�5�}�t�ё�F�]	
~ao.\C�k�Eg����0˞����Ti�^�Ax�`Vk���|��܍w�S}��T��̪mMUt��!.���9fj�}�Y�PX�)��s���}H]�˖��1ҙt&H��I����8�����|I]��ם�y��獶���_�(�X�0\[�^"�z�9��IM� I0���ԏ4tv�l�ν�s��U;46��R��O+'�tL�UF�ՁS�Ut�\�|��������2���tԷ���t���3D�� <@��fG�H�*x�߀�q��Nʉ�(Q��;��b�=��|�L�@N|��|(F9%2�8����Ѐ;��i2n_��s�I�A螗�L�͛L�_�n�To�[��Oy�,rw�&�z<a��N� �#{W��:�?"�����JﾥI��ǌ~n`��R�	iT�O����/�k&������&�4z�dט�w������Gl�N~)�jA( ����_�h3��{I��Z��H1c�f���2�خa�>����n8���ٳ��溂�ZI8'��@I��'��q�2�_:��p\I��� ±�sR�{F3�_� ���p� Z���I��'����0i������;�qW�;ۂ��IÙ=�H��M���8 �i��)#bB��G�_��V��6������L~���C�4j�q] ����)_��5�Y�w����K�@��|	0������v��I��RhF��G����FX�,4�?n�=���W�s~��y�.l�8I5�%�l�{�a�I�.��S�[U�JP.D���]�Tk)������7A�SWb��T�Q5�B�Y͘�͉�I����D��õ��Kht-���3Ve�=�k����v��'��Yf�Nd+l�Yҽ֗��)��������Z��e��I��CqZ��v�7
�7��K���I�5����`K��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xǩ"�4s2nQ�rVwp齰� ͌4s+�ny�T(#�I�I))����A�m�(1#��Z�����XP��ȭb��v݋N�����Yգq����%��/q|��]��0�ȍ�x�>c��w��'o��b9�����)^s{����иܖ����S���0i���R�&H�����̜�I0���ԏ�.fOe	��f�QaK�P�y� "X�<p�Qd����uXӦ��9���I5�4`UV#-�[ҭ���~����'n�^0o��N:�@?u�hk��Y��A�m�(�֟">�#��"5�o٥��e���\$���<3�zE�-~}���%��/q|��M����A�m�(X@�9斻	zL͊�q���Z����p��R�}vJ^ �5�h���.��&GZ>.�0S'� �ު���g8��� ӫ/��m�a��ya�X�Aj����U)+N���Ix���Ka�R8�ܻ��\�vś��Z1`�N�ǁ�f�T�B����$Ů���zւ���MȜ,��Sq'��kA&4,� ���3�ҺIÙ=�H�8�>r&���R�}vJ^�k��76�Z�u2ۅc�t\�<��C娤l����pQ/7j�F��2JHn��z�C����f�SG㴊�?����q5�n��۷I��L}JB�1:���0_hW�D$2���7 E�B��uѯ�O�x z�Jm]A�/���s��m�z����9C��,ў1�ˏ�~ǹ�z��hbvk~�#x��%��#��#���F��-��j��͌4s+�ny���.�R4������˫p}�񥒐&d�X0��A( ����_�s꘤�I��-�3��&Oa9Y֪{���ɖ?��_T���a�aq�������9X�.ᬵy��j��G#���%��/q|z��V&m�����'�>z�/^;؊��yɁ�U�4];ˍH�N"�l�V�����1�so��d�a�e�����c��%$Z'RpW��eB�1VV�zcj[�?�4��ic�v�QZ�?��
���O��5�ϟvзq8�Ј؅��FJ��v%a��!)�����f�ƳaBA�u����`�1�aw����̬��z<����]��#�z2�ŕ�+��/؞�{��^:���KH��˂�%(@/^;؊���)pL��1x�]�V����ߞ�K� �0��k{.Dt�0�Fc�<5�s z�����˫p}�񥒐V�zcj[�h�]h�V�jsUD������]��#�+�9R�зq8�Ј؅��FJ��v%a��!)�����f�ƳaBA�u����`���?ͮ����P�y��3� `A��~E��=��*87���l��P^���֮���"xC��-�T(u	M^�.�/�92JHn��z���7帘��3�=r����0�i/ȇ3
�v�v-}�	mpŴY����;���NA��sm.�9I��'���p�+m*��"Ϩ+`�|��K�z-/����IÙ=�H2�LpOJEl��Q�P�]zm?9ۄ��d1$�Q�<om��7�4����5
iEE�Gg�{�]4�W/S��8(�E���Kt�+Yi=��o�IÙ=�H�R���w(��ES���v�8:��|`��'J�	�LÆ��E� )�&�2���O�}��M�+�'�̗�����L6)�Ey������i�s̍�(��g�{�]4�W/S��8(�E���Kt�4O���x�1��&vl�JHn��z��p�Sg�3�z��SR:g()��ikp���H����Q#�?���;���N%�:+W���݇4�a�Ȃ�u�.�1�a-���7a
��r����~v���b9���eSܥOH�&q^�`
�c��><�$�;m#%�S���RY��.ZVRѿUJ��\���^�W+`�x�oP��@t�&�e�5
�`#_G����q�41&q^�`
�c��><�$��;mQ��8���/�>�W�Y��G��x�&+8@V����L��\�E�V�6IWJE�r���秹�3I^�v�%j����L�de��-@��F~*7���&�_���/���l���F�8���/����RY��k�:A�	S�r��AR1<�N�؆�B��W+`�x�o���{��&�e�5
��Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX�����/��&����H���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8����ٺ?�R�^Ƒ����"X��[7��Eb�qz�^vh;:��B�5{��
��D&e�2l��4�y��ɦ�k�:A�	S�r��AR1<I�0�f�#�Օ��qvdЧ^{�j�g��U-�e��`�?��L��l�%���V���3{��m��rr��AR1<�N�؆�B��W+`�x�oP��@t��4�u>ο��D��$t�գpP�l�L��M�,���	N^�U��ߋ��@�$��Xo��GR��)~s�����j�|��IÙ=�Hw¹��<d�7�
XǺ��g�,P�n!K��tf��
_�n�@/%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��ct�:��RE�QS����>��"X��[9R�A�m���(������{�VwtZ�+�������I?�"Ƈ5����`Ke,fi�U�ž�'�t_�GZEh5���'n�^0o�hŁw:����v�8:��|`��'J�	�LÆ�c�9ʼ��$�G�nJ `1	�<�����!�F<�+P���I��ž�'�t_�B�uʡ p�m~|��;~7����WF�r�f�t+Yi=��o�IÙ=�H��w�K��b�����(`��ү/�O'�=�eX�
\;�M +�gf���a\Y���c_����+#��.X���*"v%)��Qcm hP"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y���Ӻ��C
�y�yi
Y�2}�<��b;�B�W@:`D�h�#�*"v%)��2������1��5�;-;*�7��\@�iz��nVub]߹jGy�ˆn��?g��s>�=�+\{Yh��|����=%+]Bo�A;h�F��O�i��Ե�"xC��:��]<}J���K;�{�&��Y=�ĵ�"xC��}Vq$GѲۯzD[�'n�^0o**�ХM
�?�p�5��9&q^�`
�c��><�$\@�iz��nVub]߹jGy�ˆn��'5 �{B6$��O�&��;�L���9�D_�3���U_�+X��?<�����z��d>3EKrM3�V��g
*C�c�.[K��m w�wAk�Ya�����&��Y=�ĵ�"xC��-�T(u	M^yM��5a�)��\�v�g�W�I�H�¦ʹ
�֕v�՗ɕ�a\Y����+���LQ�X�E��uky�ѱ.��tGy�ˆn����N��+�j|j6� �T˳͠m�xW��-#��klJ�V�Gy�ˆn����N��+����]��/��=6�s���"[��g�7���ìT�T�D��ao.\C�kWUk/y@)�'n�^0o**�ХM
����@tD ӫ/��mR�MP��G��E�hxǉ �Ş(�/�K^b�Mc��_�j��i}q�^r�m�����ч��Z�Bh��vJ*�Rs�08�b(��[Nێ>�d�|Z�j��?�N�@E�Vm�.����O�<om��*)�)q	�cY�~�"���ʷ�J�	�LÆ���#��5q�ЀY@ɓ�M����*��1�G�p�Pv�?Rr�f���,(���B���̴_��EI?�R��n��am�Za(􆿳��1�Q�/L�9d������K)zum��3A�)Oqy�&�CA�o�R�GI$��ǂcY�~�s<��MR�vH9��!e�<�:ӫ���m����������p�m~|��8yL2�����ތ�1��\�vŶ�T���Ĉ��r�]@s��I�λT�v��1���2���I��'�f�Nd+l��_]���T��\�vś��Z1`�x�y�Zglё�H�a)ߤ/؞�{��U\��,�v��|O�\�+�q�� 6x�@1#��Z�����XP���f�Nd+l5����F���
�v�fp�m~|�֚?��]t���Ʊ�_�eD�I�1#��Z�����XP���#���1���Q��ǺΕ�|7J���U�
wl�G[@���j|Z�a�P�Fpwe�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL숬W@P͊Y�7#�xI��;mQ��8���/���>k��HB8�	Sc׿Z��A�.ݵ��]}�����ǩJ�9~0X�,4�?n˩�Ϊ����+p[a��*��O�t�L\ ү���f�qNS3�I��'���?"3�m�����h�n*��(�1#��Z�����XP���SG㴊�?����q5�n����a�-�I))����A�m�(Qce��ȢF:����Į��KH ���"���e�S&|���BY��l��=5;N�����O�%��/q|O{��%R�A|�stUy��DbY}n��^[_�e��IÙ=�H��=!ߎ�΂l��=5;$]��Af��s �%��<��x�>c��w��'o�c�.�09m�����
��\�H��/Sg�w��'o�V���"�V���Q�9eY��b��(�F��`JHn��z�V~�#d�	���}�pIɽ�Jz_���0�m��Ϥ/؞�{��ޝ
������U��R�~1#��Z�����XP���K�|q��=H��6�����рӚx��~ ������D>QJ A/��g�đ\e�y��3g��y����Z�� P��\�v��\aьIR=A�;�֋`NǙ#Y\��?�l~�U�{}��*���M!󂋷�(����C4'n��=?���͞��>(�J5l�����+���Zz*��5����`K���}0x��F�ԟ���Gy?�p����=R%�Kw	�F[>�y��W�}�|3����"��q�p�m~|����U0����d5�:�w�+���LQ��U�"����92<ZW`���<d���;����������r��E1�;�>�t$nXZh��\���'����%�a����ǕGF��a�1�Z���=�Ln��S�W�7����KPy]/�qF��G��Q���'��{ �=�%�*�]�1ꘐ�݇4�ae_�d
���ݪ��1#��Z�����XP��ȗd�uY��K��T��p��`�Q;?�͆�%l9�e\EV	����w1�'l�%��>/Q١Ӿ�$d��I��f�:*��v��o̙HxҀ9�@3��}th��.)rL!��di+9DjuU����Uxc���ł\�ԫAJ�T�q?�R��nścp�B��ҍ���������zP�����1#��Z�����XP������0/�e��9�S��8�U]k�(���B����_T���a�aq���U�n;p�m~|�֙X�D��U9����u�I���'����=���a���œ�,���%�a��Ϊ/�^�`0M�/�s���'n�^0o߲�}�{�%��/q|;��c���X�����w�JHn��z��S3W�K@8`+*��A��}Å�S�9o��*�w�+���LQ��J'�!�����qԏV���"�V(�b�|�5�ȧ��i�}��ڻ1�O���-�SIÙ=�H&I�3�b�}�IUr��Ӈih�|���he��G��֥��ع��&j	Z��pDY~��G��5�j�B���� ����H�ʱˡ����V�Ů���z�X�D��g�S�<�c�V�f�;���'n�^0or�.@,j#-�����1�����.��4�F1����������kר�'"I������Q�2i��e�����H����8�N����<�js��0<�%��/q|�-�(���$3 ����.`�$�4zL͊�q����1�9�\I%ji�7��
#>:��� �rmd�&l�����H���sJ*�Rs�08�b(���os0c��ZLN�	��2�V�a��h �x�����p����wя�JHn��z���7帘�f,�s��Zrt�\0�{�ms�A���S\�H��/Sg�w��'o����v�]�Uʚ7�ܩ�.fOe	��|�T������~RK܃��hbvk~�#xeayA���r�&U������G|M��'N�KR���c&;g���!a�`:O���1#��Z�����XP���B�m�/gV�gK����1�*S�b��v݋N������oV��'wNF:����Į��KH ��*PX�KL7��Ѹ��R["��J*�Rs�08�b(���zY�l��R�}vJ^�?�1�{{L	�0t�VW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�pl� �PP��ƿ�c �B�dH�7DR�i�Ρ��˧T������X�p0�&�����Q�a5���nXZjwi�U���Mչ�����Y��n�Z(Ρ����u�PBxN��X*d��Uf�Y9��_QzMy㥁�hK�'�njVfV)~�`V%'�\�*�c�-@�dƟ�&7��"=��Nc�&�Ia�΁�a�n��!�`�(i3�n`5�fK��@5���<ZJ�hEc�>���gZsT)!�`�(i3!�`�(i3�n`5�fK��0z�cUL(���r�<Uee�N��������=��*h}Nw����
�t�J8I,t�A9�AD�of�7���A3�(N��㎏qló��@d�������e!M^С$���v�|[��5�e`��9�����_�t�y�p[���d�٣���������ݹ�0�����7=����2PW�uD}%V�����F˯�+)�F�������T�\ ��i3�|)sՀ�23
������?�`d�ƇBHx\�'���Xw s4S�'�i��`�z��Y��)�?Z�����1�����NR�^Ƒ����"X��[��Q[R�75�e`��9��əS\��O�=�Q���d�٣���������ݹ�0���f�Nd+l�Yҽ֗�?��}�ͭ��I7��-5��6��	���`y���pzl��a�a���k�_�aY��|�p�6��Hh�]�!��M8���	D%��_�ͅ��I4��欱���j����B�:|l���������CyW�f�tR�wX��J�W��7/�2��2,��g�ܧ*y�E����F!K��tf��
_�n�@/%{�;����f�kN�ı��U��+�Xa�H(�˕-+��B�G����n9�}������ݼ��s�G�7s�9���on�-�6��
�jW��D���M���o�G�m�?%^�����I7��-5r�p =(�a(􆿳�ټ*w2�56ݓ��E���vj��$L�>��07s�9���on�-�6��
�jW��D���M���o�G�m�?�{|*�"�Vx�%L��W��_�ړ8���/����,DTc�~y��i���n���gW���D��g����H���	N^�U{xN��i>r�<Uee���R�}vJ^�k��76�a'�<� \�� |+vܽ�Ϝ��*@&���+�J��Y�{'%s���'���ը��_�\G��4�	B45ƃ
ᾆ�x�T�\ ���|.�Tӏ�푧)��������Ē�LwʅK�'���Xw�j�7�����0/�e��9�S'6���;8=�g��U-�ez�r�6�<n��nN�6�ϟ��n`5�fK��0z�cUL�8� �,�����°������R�wX��}�
�?�r��gGr�`@��q�'���Xw���,D�Z5���l��Vm]�]�!��8�$LQ����ɷ���/s�1��p"�,�>E��P"G�wk�١��	;q�J�� m�h�5,Wlr�r%)cA�z���a�R�wX����K�Q�4br��yO{��`�
q��T�ٮ|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/�a'�<� \f���ѩj�Q%I4���kN�����~\[$Q��
�`�ю龤9>(�vgH����8�Ј�&��g3�g��U-�e,%�0g��Յ�HN9�VTҝD!u�E����FAԢ�a\��F�dH�Dj���G�Օ��qvdЧ^{�j����#oM������ݓ��E�S���%��ì�u"4�E��b8�"e�<�:�t8:���M#�&���Z02t��S�D�����X���*"��Z�w�l#���i�ɷ���w�kkr��$X� .�/��`~�ߪ ��e��R��!kr�]Q�I����y�搲)���$:N�8.����6�Y�r�7"�p+�@���5���u�L�xZ��j�
�iB{�Z�_�+��tI�F�;���Nk��}�y:�8���/�a'�<� \�;�m�PV|1�#��d_hs�^Ξ�N�@E�Vm�.����O�<om����`��Cg�j*8a�.&�}�z73���߈�90�z��d>"I�`�c{�.ᬵy����5�t�׭��K�Q��萬�]Yݼ��4cGy�ˆn����2�-���J*�Rs�0�5�N�~u=�����z�Hi�����J���e͉�Xk�b��v݋N�����5}	��D&�}�
�?�����}�)r����'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,D�=P��[��1�U���]�!��	Ǹ�y85��L�@��f����k��$A�h��+Fen����9��0|~�LL�a(􆿳���2����.\�#$�ÙA�B�r���n`5�fK�\w��0]7��"=����B*�9u6�|�fF�AԢ�a\�y�T�g}�Ӄ�Q[R�75�e`��9G$�ء���Q]� _ό���.�}�
�?�ʬw�S��зq8�Ј'���Xw���,DH�v�����] 1�0µ�]�!����w�Հ�*��9W��}�bo{W7s�9���o>��l%i�-ݓ��E���p��b����b�g�Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/���T�/ʍ��)�`E5Xy+�Mk!P����!�`�(i3xZ��j�
����d�R�wX���7�b���������j𛚆z�Ji��U,�(�)8���0y�	�z��SR:g()��ikp���H���F`���G���`y��������5O�KlAP}k�`�B7d��U,�(�)8�}�Y�ןw�8���/�<F� ���Ձ��H��?��m��M�h{;��Tb���/؞�{��No�JH]���oAB�E����F}�=Ll�����&}0�@V���"�Vh�j _ש���yb5���[b�I���Ψ��F�wc�}�![B�
���}h�[�u O	KA��߇5����`K���ػ�T�p~z�r,J����!_�IÙ=�H�8��6�O���it	�Tߦ^Cg��)1�q�ܲ�xΠ��yGb�dW���bhbvk~�#xnůc��o@h�5,Wlr�r%)cA�-��h�m ӫ/��m��?�4D+w�����������f�l��=5;���wGu�ܝ�s2����˨(�V�֪��o�� �}��2m���l������L��@X�hD��$_s����z2�v�~�g��27�*Y=���į�4 _;��i�1@�f=H5H�n��cM�r�z�IF�˞�Bxη�H��:�-).^QQe���b�q��T�ٮ|�,
���h���J	�0�ȷS�J����Xa(􆿳����d/h�5�G�GY�)�}��EXs70��lJ��튝�b�Bϱ���w�K�	�<���BSG�p�P��<jV���\�H��/Sg�w��'o�6��T���7�8���/��Y�r�7"����#!f��$��
�5L��m}I� �-5$�sD$��y�,��1��'�al��p��g��k��i�l����@����gG1N����F�m�^�r�Ϊ�?��(��I@1���t$I+��f�kN�ı*�7`����M�Z���	4����/����DP֞ �X�m��{�Kd#���x;*�}Ւ�~ܔp�l
d��U�9�r�<Uee�N��������=��*pzl��a�)�O�=�}���N|�H�eA ��	�.l�L��M�,���	N^�U�}�g7�}�ξ���I��RhF���9���x��a'�<� \��y��`��0Exz҈��E�5��
��D&e�2l��4(�de�QV踫g(�r�N�ǁ�f�T��p_U
#W���g
����DzL㡉�&�@�}7�q��J��v1a{J��Ǻ CN��a\Y������ԻV8�I��RhF��j���W����T�\ ���|.�Tӏ~�L���vi��N�Na����g�,0 �����r�&Ɓ>i[�ͧ�?Y�Q��ǺΕ�A�m�(�hU_��_��`y���pzl��a�	�_��:�����C��֑xGV�^ɡ|z3�{.ZVRѿUJJ��.U��۩I4��欱���j����L;Л��������
�CӞD��gn�=4�D-'��7�q����d�`��	Q��[�$��X�H
$������Y��)�k������a(􆿳���Qs��������DzL�-��;���iA'R�	���i�(r]m��p�ռ�[�$��X�՚��l��H�/�n>�.-,��Sq'��_�H����K�Q� ׻�1��k]m�����9��|����⾘���c�SD釛-���>T�=�	o #���}�pIɽ�Jz_��|.�Tӏ���\42U|u='�c�-��;���֤���n�V ��a�'���Xw�j�7������7���{r���x�] %� /s��EB�w���%���ց���=�g��U-�e5��e6²]�N��&�#�(�>^�l�'s{	�h�v1a{J��Y��V�AԢ�a\�D�����R�`�|��K�z�
��vK���p�+m*��"Ϩ+`�|��K�z�Q��Y����Qs��������DzL�C��(3���-��w��k]m��F��w�6$�Gy�ˆn����N��+���o�u��"����DzL�C��(3��7�q��J��v1a{J�֋��DO��'���Xw�j�7������7���{r���x�] %� /s��EB�w���%���ց���=�g��U-�e5��e6²]�N��&�#�(�>^�l��e�eV�F��zF�ۗ���4@{A�L�de��-@��F~*7���&�__y�� ��j �0tw�*AI���J�V�	l��T�\ ���|.�Tӏ���\42U|u='�c�a����gW��_K��� X���/�K^b��6&��^�<��J���_]�N��&���3�L����e�eV�M�z$��P�;�G'Ǔ���"xC��}Vq$GѲ��W��mTS{lGD�V�B���q5�n-�@�4ڧ��~��r�pzl��a�	�_��:�����C��֑xGV�eU���("�,�+rr�N�@E�V����P3���2��:�kŔ=�	o #���}�pIɽ�Jz_��|.�Tӏ~�L���vi��N�Na����g�6���Q,|p��<_^H�z��d>3EKrM3�Vy�oY�E@���Rpy2:�׹��t��`�J9�S��˰v���K�Q�3R�e��ł)w���m�±��m|J�}�֖�gH.��2}�<��bl���>s�q?H^��2y�搲)���$:N�8.����6��J���_�Oi9L�:�k]m��,�۞��	���/y��g�'b�t	�U���C��O]r�<Uee���R�}vJ^����`a��R<�����á�~O��L;Л��|#9���b!��u��Ɔ �����Vd��[�l\�`�|��K�z��@d��ץr�&U������G|M���t�2���*!��kѶ���� ㏞ �ب*6��X#���=0Q�9oÖ�"Hi$|��ڵ�)���ͦ��^`��dg�M�q�9�}P�uB�b�#t����n>�YR��j�DI߃��K�+���w���QȘ�d�o/�d��7���ìJ���m����g/��`��ٞ�R̕q���id I�pzl��a�N��	�Ȓ�cЉ�MOc�����2}�<��b;�B�W@(��T�[�=�5x��j|�>�OU��9��]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e5��e6²�T:���V�����,Ǣ� ��^�:Z鎬�������(���`$�P.eE���lC��U�T�\ ���|.�TӏU�m#j[W, +$IA ͒�ښ�l�L��M�,���	N^�U{xN��i>�/�n>�.-,��Sq'��_�H����K�QR�Xe�������(2���􇃬Tk��A3�(N��㎏qló2u?r���Y�G�˱�ߓC娤l���Mq&���[�=�5x��M��%LS�8o�f���k�:A�	S�r��AR1<]Q�I����y�搲)���$:N�8.����6a'�<� \|���yB�+�kv޶Gl��C*�󅒣$���:�kw�j��,�0�@vV��
��D&e�2l��4��a��se�`��ٞ�R̕q���id I�|��{>��e�t�b���6U(�<"s����&=�rs�i��O3JT�!I�T�\ ���|.�Tӏe�t�b���6U(�<"�%�2C��rs�i��O3JT�!I�T�\ ���|.�Tӏ ���v�l.�
��ڋ��Q]� _�rs�i�CЎ�����Ɛg)x�D�����X��Q��Y����Qs������T�e�V0�� ��vзq8�Ј'���Xw�j�7��	3i�\��׹��t�M��|S�/����Øf��K�Q��`�����!�`�(i3�d�٣�����6>��JX-�ܶ�0����K�� ��^�:Z鎬����Y�V��#qX�9y��"Y����8eZ鎬�������(���SG㴊�?����q5�n�@qQ�ܩ�8���/�a'�<� \纅<S�O؏����:aޗ�U$�'���Xw�j�7��	3i�\��׹��t�M��|S�/������������bpO؏����:.Ɓ�dd?QZ鎬����Y�V��#qe�t�b����t]������ī��]�!���1����mA<�}	��G��[�f�]n�"��V��d�٣��c�A�L'J����l�!��G��+�c#K�e m8�8���/�a'�<� \<F��̎ÆLx�A�B�m@�:\*�Z鎬�������(������aU�����w��T�\ ���|.�Tӏ�'�ŀP��3B�\G��ﱴ=�]�!��	Ǹ�y85��5m*�Y��g�S�<�c�!���X��`y���pzl��a�D���ƨ��u��u���� ��)p'���Xwa'�<� \f���5���w_������8T��]�!��i��&�J@{L�'x�$vcH���K�Q��2�����z��I/r���+b�a�&!9�q5 ̬����b9����Z[Zz�! HڜԎ���J@{L�'x�$vcH���2�1L+�&!9�q5 ̬���M�8��;[�(��Jx��'�!�Ѣ$X�jl�N� �$]2�/.ePN6����(�;UW���g��'�|v*�n�6��.���I��N�\Ӽ�gy�A=D�!v�w�u��.tƙ��3Ve�;�0�XǷ
�J8����d��MT�D�9�.g^�F���p>�����;mG�����k�}�m
ˈ��$����q���w*��	�a��������t��P�mjS�z�9U�s�Z{�=����X��-��sޛԪpP���4�?CZ=x 
~�F�踫g(�r�N�ǁ�f�T��p_U
#;��|B��>>0j��Ih�	�;��J�����M���R��ӟ-�F���ˏ��Z��zf	�$NT�I���I���C1zh=E�g�N�������S�_
�u��Yx�I���I���C1zh�6���Q,|�rHYSڣ��ǡ�C�a\Y����+���LQ�s�xV��8���&�@�}7�q��J��v1a{J�?��кDO�,\���ӟ�X���&�@�}7�q��J��v1a{J�d�	@f�u �U�N;k��!a�tc�&ck���>#qBK"6j�"Hs���ٚj�ώ ���]q��J��56�f�s�G��J�����M���R��ӟ-���4�&����Z��zf	�$NT�I���I���C1zh=E�g�N�8�dEm7�w�kkr�I�;(�\��8p���uAԢ�a\�DW��E��q�����C��֑xGV�eU���(�CK{D�sss2����`�|��K�z˦9��iժG�p�P���ً ��3R�e��Ӵ�"�6j��;٬sf.�5^����r���zk2�����n�۴�.�<Mm1���P�|T����E�E��3�L����e�eV�M�z$��P�Ġy�����l�p�H1�a-���7a
��r�$Dc~4�A)�V��/�c����sL]~цt�U(i��[���P��d��MT����k!Tޙ�ǗL��	��q�©�����<�������~s���^�����g��,\ަ�It��+g[�b�ӝ5�T�w�%b��Gv����Y���a\Y����+���LQ�~�#UJh�������\����>'���������6%�a�ٙ���O�#t%zY#G�!sH�\�t���\�W�D��t�!z�t�-$�I����Q��K��::A9�C���=�Ҹn1��Et�!z�t)P�a[)9b�jT�.���I�]�Bb���{��¸�m�B��d���m l�o�@`�~�&E4@Q�/�9��?xsl��)��'���Xw�j�7���3R�e��ł)w���m�±��m|�vA�S����A�����~W��� �A�J�e�!�c�A�L'ӸT�?��i��N�Na����g=E�g�N�;�/B��[b�0<��U�%
�b~�1�W�~�`�S��P����{�j%a}�C}��0Ex��L�.��W��2�H=�m<����6U(�<"�CK{D�s���?�Tl���FѱTW%#3?���*��u�Z�	9]�l����l�� �qe��E��'Z*)�?�R��n��h
:h����t�h�x�܀�>5���c�v�_����J����/g~�
�97��ENҽ��O�ʦ
���c�v�_����J�����&����˶p�0u�xs�&q^�`
�c��><�$jI���RUyX�C������u���'b�'=�(8�����FiŞ�W�%3AԢ�a\�DW��E��q��u���'b�'=�(J�}�֖���J�_��e����7���{r���i���A�@[�_zβr��o��SO�W,�P Or��mR4���oP� �qe��E��'Z*)�?�R��nj��P_Q����t�h�x�܀�>5���c�v�_����J����/g~�
��C�|J3J���\&<����29��#���,\���ӟ�X���&�@�}�-��w��k]m��+qO1U�)�#qp���W/S��8(�E���Kt�4O���x(��&/�j��8=��2��3�L����e�eV��iA'R�	.s�b��O�4br��>G9���ļ���/���b�Bϱ��3R�e��Ӵ�"�6j��;٬sf.�r� F�3N����Od-@��F~*7���&�_5�NS�x�r�r%)cAS�B+����;��|B�����
:��H����_��v~��S�?�o�ߚ��x���'HY-��Yk"1/s�\"�����p"�+ڍ�P��Gg���/�9��������֢&@��&;-;*�7��vє�&�������7���{r��W�Ty��5�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��sI�$����G[�� ��aP��k�= ��j��C��[�����p��@L��X]��U��|5�.4���Q��K��::A9�C���=�Ҹn1��E�<��R�������7'7�}M,�d�}}wS�7�}h���	;h�)�[���6�5�9�(���u٪��}���t��˳�M[�����'B�ɏ��]�!��	Ǹ�y85�0+ע 5N�I���I���C1zh���\v2:R�*��&��K�\7}�W,g�%Y��̗0z�cULj� 1ɡ��&�@�}7�q��J��v1a{J�Ӕ���(�q�\E��0�-��*�6[�j|�>�O�|���9{k�h�+�d�)bU����,ǢL�E��<U�����9�4]:C�2Y~�O&�r�$��3~�����2V�a0��r�N��(�����Q}mҁ�t����s}�e���dz�r�^d���#S��d�Q_�;!��i�W���3R�7�z��?l?�d���&�o�,·��4����z��kɡ�ܬUvd��� �D��$��p�����"e01�"V�����a��"�qg���0vE�So����~�y;z��y7��8)b����ߏ�U�ڴ#�������g�+�è�P�/7e �v2R�=4�a�4�ĂB
S4ɰ/]i�G��'(�wy �v�0�*'���C@(�tW�
v�er�� Wl��5�9�Z�8 gV�A���r!B�b��T�Q5{d���壟2$6�sIEk����V�a�I�.z�[o�0_���E��)CI(�0 ��,ה�u�j��U�T�#���	R�%�MK4/�[ʙ{�+j�!����$\ �h�q&.&οiboI���Hc���o����I�AV�u��0ݷˣ%#~��m �#g�k��������e&os�@����A$�P������5d�=k�Rm��̬��U�u!�?8��Cd[U�8�h�DI�����[mߍ�C*���M����{_8�Y��=�}�Vݨ��\9�oA�
��߼L�T��~��Uг�|<������M�h�ˁs��Qf�A�������[mߍ�C*���M���)�O�=�}���N|�H�e�8�m
��NjX�U�4�04�jf�5ߧE4��Fi��|��6](���T"��D�t�$+���t¹��R�[vf�t��g��;X�-�!����~�d+[.!�ώ ���]qP��1cdh�5,Wlr�r%)cAQ17�b����#g�k��K�c�\p�q����#@�Q¢�r}l��L��M����,\���ӟ�X���&�@�}�-��w��k]m��+qO1U�)�#qp���W/S��8(�E���Kt�n ~���7�� ׻�1��k]m�����9��|0�rI�yV?�����P�|T����E�E��3�L����e�eV�M�z$��P�^�6�V���Wy޶�W/S��8(�E���Kt㲓c�X0�jqV��	��y>��
6��Ih�	�;O�=jʙ�4�-���G$�2����� ���JH����8����F)�~����H�V��^�5G��-��;���iA'R�	���i�(r]��0�|����񔖔�c�fi�d>G9���ļ���/���b�Bϱ��3R�e��ł)w���m�±��m|J�}�֖���J�_��e����7���{r��f���꜅�R��ӟ-�|qU?R�f\����Ô��v1a{J�w��7�ZEA�U
/c���us\�o=S���%��݈c��ʨ���z��F}���V6��Q��&i��N�Na����g�6���Q,|6Z`8&߅=�(3�Y�4�&q^�`
�c��><�$("�P��_��3�.�J�|�+��?�d���&��$ͯ���'^�!�m�фX;<Pȣ0o
zVcP��CX�|��x�^:����3�k�~�f��*K��P��op����=}'t<��ġ��,�B��(�=�g()��ikp���H���3soo�ۇ^���\�}w��7�ZEA��&rm�\�K>e����m��+���J q�v����6��w�1���|��٧�\�T,b0V�u�Qi�FkmG'w��á�~O���-@t�/�W/S��8(�E���Kt�8�T��fNߨ+����qJi�];���w¹��<d�J�^�l��?�z[X%�88�;矷p�]3t���m����5�}�]������2���񥦢$'5�J�~���.����7���E���b�jT�.��(���m�|b w��,�9)��j)yc�n�.�_�t���L57��DgR� �ұ�X;p`�gR� �ұ/EI���ā4@Q�/�z��1$_o�l��)��'���Xw�j�7��6��~p�=�J����6x�F�-LU����{����8B���z�!��ސ�n�|����Y�{'%s���F�\����Ô��v1a{J�w��7�ZEA�U
/c������󾑸&'Ƶ�s�-��*�6[�j|�>�O&n'o��W�N��x�����	p)�O�=�}ҝ]��w]3�����������V&Fndq��c��	���}�:�>�f�T�Ĳ�)Q�XI��J�)���3J�~{�ڲm>>*�����*[UxG�#�9�[Їa�/!O���锴�;��|B����j�ݷ���1K�Y�bm--��'��m�*p�<��y�c)�h�<om���Z�,�h(N��"~6���aq�����!�G���Z�ה�	��ُ9l��w���]'\gWg��	�Z�kfc�Q�bc�+�(��?c�0&ڝ���M_�mS8<�n���ƻ��g��n%�)eUȯ�����J�^�K7͍��|��W&":&����1�^��C�/�nu4Bޗ��jw�	���K:+>X[�QB���X��WG ��'Ƶ�s����,Ǣ&n'o��Wt0Vo��X�m��{��$E������V)C�J�1���K���L���4�04�jfFi��|��4��U�����I�c�����M�~���y�=:�����ˋ3��=TaN�:+_��'5�?�°q�>�I���� hTc44�.�K=�^#'�������L�t��n#�%��>�r�.�kR��awfՀ���di���t��Pаe�E�k�\D!�g��9cbX�8�SJk韸�b���M����A�m�(��D׉��h�#g�k����awf�#�%��>�h0Z�W��2N!�y{+��0ExM��"f�t��b����^�;��|Bu>ؾi��H*H:Еz�=癍D��`+�CU�M*�7`����M�Z���	qb	��G��-������X�m��{��$E�������_g�$�����[m�ɲ�cz���Ps_*�GqW�w��fD!�FPFi����B�#;��|B�¸A���iJ���S�NNN�� �aw���U���p7�<��;�B�~�{�Jt��K�����	�jo�����m���m�K���/���ȜR���?�d���&�^�n��Uh~�1�W���h*
��#����[m��3R�e�����v��a�^�n��Uhql�d_b�����r�)�O�=�}���N|�H�e�{����3@[�_zβrB�ek�5W�|r����H�Z��D��!��mku�mۭ1���P"d�7�4��~k��D9�$n�,L�N��3jd��O�/y�y���"b��g��i��?�-�>�h%�"���k����K/����8'��ģ/͖��$���xW��*.埲�Uq��Tѐ��rgS��R-�iBPd��8Pb�zc0�]F:����Į��KH ���{Mý�uD�%WJo��_�n�To�[�C��-����]��������|I�ۏ^��d�;��|B<Ww�do �X�m��{�b���L�>j%J���E[z�taS��R�Xe����b�A��d8r��?x5V��	��y��I�A���U2�h=cy\��9:��	���%�� U2�h=c�ac��,����]��0�ȍ�x�>c��w��'o�!b)�C���T�T�D��ao.\C�kRşe��J�Ld�r:ha3B��*w��z�Rɏ��Z����1��]%�@�γ�t�`~��5�#y:�}"Oa/�)(�&��^S��ȭ���$P��G�T?s��������T�%n�"#( ��PF�yi�����8���%%��jr�>,���6P�x�Z Y�O`��[��ȡ�m�qةF2dv����YX�bϒd����ZkZ�y/A�T��剠X� /������i=����C�/��z0c�.[K��m㳆�����{�E�:_�˨ʿ��w���f�C�w=ء	���!4�.�>b�!H ;�|㡼�V�}Z9L�*��.��Ӑ��>��dWa�X�w�.ᬵy��(��8�\�W�w��fD*h���}�f������C;��E5��d;��|Bᜮo{Q��ȷ��>m��Iu�`�o�wqMYxw����S��j|�>�OY�^b�(���t��h�	�Ȟ���?{W¿pX;��|B�'	�?��[�W���j�S"�ލ?ڸ��Fp���0f<N"�<om��v��E��zq_<�>>m��S�-�kw��r|��߇(���л��e,w&�#g�k��R�Xe����ɲ�cz���v{��lw	����,Ǣ�Пe���;�L�t��ni��:_m˨9��|��7�k�ly�mDƝ��0vdLqgF���~�)V��B�1#��Q����Nm�f�X�m��{��,M]�i{@�c�}�CL���yF�� ,��rQJ�ڣ.����X:�@�7"�_�Z��E/�	�Nw�A�Md�sω�f0� �E��'Z*)�?�R��n��h
:h����t�h�x�܀�>5�[�s���J��sr�l�k]m���+}8���97��ENҽ��O�ʦ
�[�s���J��sr�l�k]m����ǡ�C�a\Y����+���LQ���ll��4�(�hF�w���a\Y���o��[^ �﵇zb��B�>��֑xGV�2��."�z���`��vAԢ�a\��?�D�p&B�>��֑xGV���KKH���&q^�`
�c��><�$N�w����H��4�d�cX~|�D́.�.����|�+��?�d���&����|��+�+\���]�5����V�f0� �E��'Z*)�?�R��nj��P_Q����t�h�x�܀�>5�[�s���J��sr�l�k]m���+}8����C�|J3J�Q%I4���H_r܅�AԢ�a\��?�D�p&��2�ę�u'b�'=�(�o<4y���W/S��8(�E���Kt�4O���x�'�������p�+m*��"Ϩ+`�|��K�z3�_�並ɲ�cz���ł)w���m�±��m|�hU�AG�����zk2���dE���;���]�F}���V6��a[a��|u='�c�-��;����W�O�힬���7���{r��f���꜅�R��ӟ-�Wڭ��h�Ɛo�c�?EcD�=1]M����_�@[�_zβr�j5�{��2��@N���#���
ɴ��z�4�	���WdM4@�GhC��BO�]�!��	Ǹ�y85��m�AD���"'��l������O2��."�z����&�@C��(3���-��w��k]m���@~��&�v'���Xw�j�7��ɲ�cz���ł)w���m�±��m|�hU�AG��.+�x:.���͉���������&ea�8��������?9�M�Ч��Dua�\����;��x�l��1:�N�*�xA�sxW�O�Ji�];���ss2����`�|��K�z�
��vK���p�+m*��"Ϩ+`�|��K�z�#$�e���w¹��<d�Ji�];���w¹��<d�,��L��T^�`T�W�88�;矷p�]3t�}i�@�5�}�]������2���񥦢$'5�J�~���.����7�*���<�Hr��r�,z_�����9ƿ���=�Ҹ��tk@�Zۙ��A�>s��Y�&�������t���c����8-�ؤ^~�X����ɲ�cz���ł)w���m�±��m|9�n�����U��R�i����C�C��(3��7�q��J��v1a{J��Q�v�(��d����==�h�f�������m"�s�lo�������	p)�O�=�}ҵaM�B��5�Jmf��4]:C�2Y�/�B@������Kb��r�N��(�����Q}mҁ�t����s���#e-��#b�^B���B[on� �I���� h�����S5Kȷ��>m��Iu�`�o�wqMYxwN�H�� �\�a�G�r�B�$�N���$����Nv_���GXE��z�Np|��T�����oȊ P�������Q5r�����#T��hT-�X�3��`�ձ�ʽ�mT3y���I�d��E�]IH[/p����x!����<�����Ȕn�NQa"_�~�c�To�
b�
jPV$y2�:4Ǒ$����NO<���*�m��Q�9�o���R���q��W!L�Qՙ-��2�O�$��ꤹ"��{���}����bNm'g�1��
�q���cŘ�/5���c��Ԡ�~\$#�[�#������W��͌Tf�����Ȕ���8���/��q28��y�[�u7*.埲��Y��"����:�5}`���&b-�.���������~x�k�/�x�˳�Qx�P�������ATm�X�4�%��^d���#Sx�z�/�Om�#��H�{\#ȕ���v��R��x2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�D�{�ը7	�1�_u�b3�ڪNTRlj�Ŗ��g���kt�Y=�R�}P,�?��Kj�^��+5$!�����6�{�5}'Y�:��w>��Y��d���!i!q��V�<L��-�Mφ�q�©���?��P>�.�z,yPM�^-q�x�l��1:�N�*�x���N�4���f�����Q�_f�Nd+l�Yҽ֗��k�+9=�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=�m�n���֣��n��ݜt���,\ͨ܉p����O,8�ݚ�Н�bs��2[������	�;�ݚ�Н�0q���Q�L��
�:qEp3?���*�YmC,igu?V��j�c<�s����	��7��u���/	�C\�2x���?V��j�c�?�#B,��	��7���=��ծœ��K����f�?ǉ�=2W���R0C7z���.��.f���T��M5��s������>��>hߵ�V��rU�w�⽒���M����A�m�(��D׉��h�#g�k��r��18�� TF��&~����ww¹��<d���lC��U�T�\ ��;��|B����=���p�� �&SfzF�.���tAC�����[m��3R�e��,z*ը����u���"6J���_��ocm����$Ȣ	!��.���� _>��>0i��.��J�������^�d�����w�>f��8�Dw]r���|�|P8}Ά�ud�H�A�m�(*��l�- ��pg^���W^G�2y���H�V���b�?C�F�.��.f�Cz瀿3�z���]�D�)�O�=�}���N|�H�ejxL��Ƅْ�k&N���g:%���5�>�k�_���(&�c����7Q{��̯Ǹ���)/04K��%�&n�i��V��yRf.ܸ���=���G����*�7`����M�Z���	(@��,1����Ѹ�Z{}t�\mc�#g�k��7�_�ܦ��X%�(�!g�lu/����t��P��M��%LS��b���jp��0�| ��p�-a�D͢?�d���&��bya�C��<^&!!HY��w���V��	��y�� �P�qN�h���w3&�4w�d��˩���.p!�'���4��Ǳ߁Ĉ��r�]@Oz)G�F�C�T�\ ��;��|B����=��F��׿]�v����D�ه4�tZz_nÑ2hꬺ��1��NjX�U�6j�"Hs?�Jy��{Q/�C�#>��G�Ȧj�E��g�Hb�t]�<Lz�����=�<��̀��unЅ����D5�|أͽgF"?f�Nd+l�Yҽ֗�,�3�YG�^���\�}GP��_&?Wcv�mAvWދ�qc:ct�:��RE��W��_��MM
��,=?�d���&�����x������v
6ڑ�I����<�W?�I��RhF��U>V%`�~��POۭ�٤.��.f�Cz瀿3�V���!�F?��G�Ȧj�rZ�0m�\�n�8�Z�Ѽ�;%4fC�6j�"Hs�2�p��΂�j�|JK
��ݚ�Н�Z��E��3?�d���&�o3F�ȧe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI��ߎ�x}�IUr��Ӱ8��oZ<8�w\�PPOi�<ՐW��K1Y-r�EHd
0Ki�|2;$�J��7�OT�,��7=����2PW�uD}qb	��G��	i5Ɨ�}�IUr���v ���\{a���k�_K�ǟ
��)@[�_zβrꢯ�wv��QX�mR�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�wP-�H1�m��d�7��dt�{��!�r��I6�qf���?v�q�2�_:��p\I��� �W�G��!?�d���&�db�\EXP-7�vqq��I�?g�f��r�F�5��I^ξ��ݴg��S�ZC%`Y��V)���n	l��Q;�im��ȍry��	^�R@Κ�2���eip���,��x�y�ZglZ�(�SڬG�ݚ�Н�3A��gd�J�`���nU�gF�r�f�t���MK�L���NK�3�Fq)~�@�&-)���(`��ү/�O'�=��k�+9=�]V�H7'�R�^Ƒ�ӭ�i�\�>&�&i��	O�^
D�5��Dz���X;p`�]���!�D�-��60eq6�oǍڍ4��Į.$�L/���?T�x~1�@����Ի��= ��j����X�u��
)\Y����i�\�f�~�ڳkԜ93�����U�6n�jD�pϓpy%����ڻ�<i���eŞuT ��>��p����nZ���t��˳3[�u8��⒍~���*IϢ���z>�6����iA'R�	�2�O
�� �ݚ�Н�+��%�k<r�`�ab8IU_h�7��m�K��ݚ�Н�0q���Q�L���/��@��e:$h�7�cl.�	�C�
�:qEp3?���*��+kt�Oz���)���s�������n�r�\E�6E�
0�)�ރ��(��9�'b�t	�U�F`8m<����վ��lb���V�G�i����SzY]�埅��!�ٞ�'�/��T;��%YM�	�v�3�x�y�Zgl,�B۸��f>x�:	�W+��W��g�9��,Yb�;�
[�&~����w��FH0M�F�r�f�t�ŝ��X��MM
��,=?�d���&���=����t/�������� �mD!g�lu/�8
l]]y�1�b�'Be��sߍTl���g��b�w�R���ykb>���p�������nSf�Ǜ|��LiVݳ���a�����o��8q��ǵc��5�%]����8�B���ow_;O
�J��:�����nސ���B�ӗ�z8
l]]y�1���"�XNAA����E�i�m}66j�"Hs�ĖYS⪞mf��aT��3G?�d���&�zY]�埅��!�ٞ"�_�-U1�.�g3ZQ�ͼ����GsG��*�7��j��0�h��7n)�26���k楊HaU$kX�.SS�Zs�c<�^<�H�W+��W���	�|Jgq�M�4�9�0��L�w�R���y+1����!���Dt��r��`�@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���ҍ�X�b�)	}�A-�����p��(�+��T��/o��إ�8p	�rh5��tE�ӻ���Z=%���X�����S���� "5�]�i�ۑ ��GZ>.�0������i�p���,���C�M$��k�+9=�p�ϵ�DE�Ʊ�_�eD�I��<P��C�Ǚ#Y\��?�l~�U�B�)'Bz�;{/�>?����n!�`�(i3�� �hҪ	n����������������i����u�UgF˯�+)�E;�G:��s=��]zŎd>&�&i�������kޮ��R�^Ƒ��f�?ǉ�=�d�uY�؃�]n������+��cy]/�qF���MK�L�t������ݪ��t����$�����p�><��d5�:�w�+���LQ�f�?ǉ�=gR� �ұ!�`�(i3�Y�M���˻��0y��<0��s���4@Q�/��y��j��k�lԇ�-{�t�%�Z?��<�ry^�h�'f R�苇��Fe#OOJd֯�|�)՜�4�X;p`�YmC,iguEOJ�uxm�3���w�@V�?ZFw�N}�IUr��ӭ�
:&��5��=����t 7�J�[�_�C�6%�W��|K:�2�O
�� �c�_������=Ro�'!#~c��n|s�)>�:��
K��>vE���2��)�2�rMX�L��|K��h���a��ƞ�{k�h�+|�c�$�t�/*;63��dn��A�v���{	��+ptA-I�p��g���^u�� 
~�F�,���XF:������X`��w{���Z���F%�X��O�_�-��0��ԡ�/$a��F˯�+)Ƒॉ,����g��U-�e a⣃_B7�}�!���:�,���P�,'",H� ��ˀч~&5�r|�g�ܧ*y�Y#	߾u}�	76�&�;��|B`#���J��M�r�!��X�.����2܌�h,\�NyVX��-|?��Vx�%Ls�N
�u�}�T�\ ��;��|Bc^���HV;ƘdO��cb>�h�D���b8IU_h�¦�naä��,bxqX�����,�ǰ��������2܌�I(�g�y��6j�"Hs�l��J�&b���J�/�߂�숓][3�X���o�u�/D�P�$��0o��]��A�ϵ{�kߗ��,�r�hr�W�u<n?E[��/xpK%����NJ�q)t�"_���I�>��t�2Pk�b���mjR}���܁���e�G�Ǆa"��<ͯ�G��R'),��`�퀁9��!���Z��L�dGk�>}�����L��Ay46�o8:4�I���c�90�Ǘa��xO.C��WHe�Q\���F�`yx�>�+X�M?��y�!�`�(i3]���!E�r &
�$JE�g�������(ӈ���m�r����̢k���"��w6�0��ɗ��zi#Y)M���Fe���2+m�7m�T��Ʈ+ˀa��z��2�,�s�Yls��8��GM��-����!�`�(i3]���!E�r &
�$J�� �X?�V޴�ik]�Ws��h�GHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�\;/4ҟ��,���Ъ�a�DP���V��	��y���"��l�����ha��nt�"_���Iw�4���x#Pk�b���mjR}���l)�_���=D���n�)�<ͯ�G��R'),��`�d��RY����Z��v�ء����Ϝ��*@&���T���dn��A�@zS�WV��	��y���"��l����:`mW��J)�h�O{2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�����o��m7n,�
��W�.��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv��T����M�@�V��l�c�jd�LdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu��"Όd)���W)�x�F[�-6�$�D	T;�i�� ӫ/��mR�MP��GX��WG ����׵���G��[�f��
�����'�^����8BW�R7���r_��m�[��l.ub��|6?����E.�`كcf;[���rw�&�z<aF�S�1 ��T����M�@�V��l 1D���M��hi�aDU�G�a�E�RD§B ����z� 'J��@�D����X�Q�j*��{�%�@�V��l����,���b�������`y����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��@qz�_vrrL�����
�>��L�?� �T�"�}LT�yo���
^���|6?������|�����X�Q����`�v�������s���B�_��:��%g
C=��Hb�8�dX�↨q�©����y,�m��M�5�� }����9e����1�:�Ω�.�&ʺr����$l����<�2^"�u��.��������֢&@��&����Kp&�@���k�֭AQ�0GȨ��_�\G��4�	B45��wxT�;�Ř�T09�����\��ą���d��Fn{�^l��R�G�)q��`^�GHN�2߄����o)�]rH����8���f��9
���M���R��ӟ-�'�0�zA�T�g�v�0�}�X~E?��#!v��;�Ř�T09�����\��%<�i�G�/���r��1�Z���=��j��6��������k�+9=	��(l��U9����u����hAI�x#2���p�����x�B0��s���4@Q�/��y��j��k�lԇ�-{�4�0 L?�p���@Z�M�g����-����b=���
�	?�<!�`�(i3���&�j�"���#?�DsQ�V�r[%�/B��亁��$-q�0c$��2��}��=�lx+~�^8�]3t��xE���8��)qD�	�	?V��j�c�[N�&ѐǂ��%D�$o��)�ͳ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���L���Ŗ6$\K��p�>&�+���LQ�����_��j��N�֞q˩���.|�YtA[���Ŗ6$\K��&b���E�vL������ur]p�+#���&�x�.E�FY��+c��8���ݔf�zE�񪣘yg�U�։�������� h9�=�^�a�	�zQ�ě��������]�9d��U>#��-䤔���8!�b#\w��o�x��o��ײ]�4�Kq%��M�Vr���J��:����;�	��o�g��}>�IM8e�׸J�q��G��m��+�Ƽ(��h�.�z,yPM�^-q�x�l��1:�N�*�x��
[N<p�U��֜��3�X;p`�Q�%�+2�j;��q,�?�Ho2��ݪ��t����$�fC` ��\�H�MPq6.����gQ'�|ݔ�3�(n�'�f�?ǉ�=$(��>��������	���i$;��|��T�.�l�.θ��q����k��,�:�N�*�x3Lv	̅���X;p`�(�����֭�h��O5�tx\s�l.�	�C�
�:qEp��:��ZL$�����:��IK��<[�л���7#���=
 �4���ߩ��ݚ�Н�p�n���d�)bU��� �Y.�.�g3Z�7�4��~��=�>�:|]η��E�<���5[�������0j|�~{b62�tstJ��:����s͟;)f���d�jO)īIX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�+��%�k<a�E�Rq���my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�6��J��c��Yu��"Όd)��;|>r:w��չ���1L��bsAOw�*Y��b"���LQ�/81tSjv��wӨj]h�jsrCm�k�`��.���'fr��B�
�:qEp�;�P�t�5fĉ>99��A0ok�׹��|�T��U�m7n,�
�t��϶C�;��|B����j��xvtL�i�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcd���;	���v�����t�{���6������]'m���G�K$xE�p4rqG7ʪ��O1�Z���=��T%O^,v�U'�W�Q�4�gX��>`���'�,A��89��A$�P������5d�������y�(����<m�r$ɓǃl[�Ƶ�1tSjv�?V��j�cF�l�q��my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�6��J��c��T	�����Va�ir�Yu�������&G!�`�(i3�$���"�U��I�,B�E?�xu�jf%���F|`�+S�p�����;���ݚ�Н�?V��j�c�:#��XB��4,�Q��U����z~��6��	���`y����ݚ�Н�$f��_Ub�F�S�1 ��H�������
q<O�A'�u������O*�������.�K{e�Il!�`�(i3�Zj���
Ĭ��,��oX��ͧ��0�u8�a%�R��6���n6�NGq�T�It���P�7� u]9�#�I�3b�������4,�Q��U����z~(ȇ%�>�L��>e0�L q��j�J^!�`�(i3q.U���oX��ͧ��0�u8�a%�R��6���n6�NGq�T�It���P�7� ������mo3b�������4,�Q��U����z~(ȇ%�>�Lg4��Qu��r��!�`�(i3�� ߌ��9f2Pih{mX�ra�R�^Ƒ����"X��[��Q[R�7!�`�(i3�����!�`�(i3�H����+�uB;y�qT��#zɯ.�]ؔVGi��ċ�!1tSjv�!�`�(i3?V��j�c X-�Y�{'%sk����w�;{�'8{1�']�JN�Zm1�Z���=������1�Z���=��n��I!�`�(i3��w�w:�!�`�(i3!�`�(i3e�v��ҵl�]�!��	Ǹ�y85����[��蛫���dU����z~Ao��m0e9�Q����0�&�����ݚ�Н�
�:qEp�;�P�t�5!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx܇1~�}��Ϙ�h����A��܆w�R���yK���}`�=��.y�!>�,��V.L3������ׄ�hNݽ!�q�
�Bk�i�����Bq��z0J�1�Z���=��T%O^,v�U'�W�Q�4�gX���^�q�g��IX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н��lTN��IdN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-j�1tSjv��H����#� �,W��5��t�����F/G��Hb� h�ҩ�?V��j�c X-�Y�{'%s��1ƵS�VX�9i�S�'�)�Բci�'�/=n��jV�{+�fbmDF�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j���_J��`U�a�(�>��(8	̜���,�ǰ6X����0敐�^p�=N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��_~�TP���V��m�̖˄��OT�<��h�l����pE\���Ja�NJN�ǁ�f�T��=JB$V�5<��D�^�3ـ1�� ���JN�ǁ�f�T��c�H �$�gm隦���W+��W��D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vci����
܇=�1h�p�i7N�_�z*K��I4��欱���j���t�0��,���d���!i[��*"�����:�#�|$.@L�`��]��8�8!�`�(i3!�`�(i3�gKh���V�H�M�[��*"�����:�#�|$.@L�`f�Nd+l�Yҽ֗��F�I7�/��gKh���V�H�M�I��)���W�w��fDl2����}*�NRcnvyw�R���yW�R�w���L�>5�C��Ҁ"���`Vk�d��f�Nd+l�Yҽ֗��Ús�Ww���M���XH {��u��]'\gWg��	�Z�kfce�E��TP�`���φ��<�6�̓@?5�e���ɯ;���{���#�0�zG�������&G�� л����M���XE�g�������(ӈ���m�r����,�u�S��d��JXl'�T��~��Uг�|<<�6�Q=y�}�6f&rG��Hb� h�ҩγpo守�u�YN
��)e���T���b�Bϱ�h�5,Wlr�r%)cA�5QN���d>�c�n�P3�K��b� h�ҩή� л��P�궊�2�����8!��?V�ы�(�)x�?{���x.�Knq'ێ����� h�ҩβ��y��lDe7g#�qa��T)�
���l�K�>�������� л�1���~!�`�(i3�}}�D�������˦G�K7͍��|��W&":�ݚ�Н�0��l!���O�D mWN<�6�Q=���F��O�ȓM�Me��&[�x�R�"�,bxqX����F��O�c�ˆ�A��߸��S�Ȍ�d�n�ͻ���~͏��a�Om�`�3ޕ ���t�T��?E-h��`f���s8����z�:Fa�7���W"�P�K¨}�n/�J� &�0D�棊�{���#�0�zG�������&G�� л�
��7t��i��nF���<�W�.�P�	��
�Q�}��b��~�F�KD�Vr[/}>5��0�B� �b�Ю� л�e<�Ia��la��o���H�RtV�^_v�9�+Ǟ�̩jv�^������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��;�uO��Bu����aGl��Z����pG�p�P�m������,���s�M@��N��$��Ɇ�����5��Dao.\C�k�2v@�q	�L�F.	-�L��&PY~�y����o)�T*�c���-/a8!�`�(i3��a�Om�%?es� e��0�U+�qbp@�!�`�(i3��Id�!�`�(i3R���Xc�
��7t��i���OLQ���M���X"���&�^��v�8:?�'����v�]��1���U�._����P�|T����{7�H����8���O�υ���YN
��)e#j�o����B� �b��!�`�(i3O��(���*�֦�n�닓.�`�3�ԝy'����y��lD&[�x�R�"��}Dq�f���Qѳ$G��A0ok��0��l!���O�D mWN��Qѳ$G�ѵ�q��]� )�+�!c�2���#Y�������0���KU�I�h��^���p����Qi�y��T6OY�=6��\l�Ud�exB#�I�i�D��%�:i>��E�N�$mg�U�ʸ�#4��_v�Յ5`�Mq�I�g�ݩOϓ�I�i��mw9���יaf��pD��A�,Z)�<��Ky|uU��U�ͪ��ڋ�9�)x�?{���x.�Knq6@Aa7KLY���F���.:���dy�}�I�Ҡ8jH�G�NJ���j�_q�φ��<�6�@a� ��`6:���ʃK�,��`��%��	��A(�c���_G��Hb,���s�Ma�"Pn��s�I���I�����OeU���(;)(F�T���L��\�vk�����k]m��Cw�Hm�̭b��v݋N������'w�T!h������)x�?{���x.�KnqO+��>���W���Ҥ��L�V�W�]=��b��~�F�KD�Vr[/}>5��0-M�O��~��?�,t�J�,l�����(4G��>����aGl��Z����pG�p�P�m��������a-6�Da
Y���@�?'���c�e�+���4.�*�l��=5;�a���8n
V~$o�u�Q��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$A�׭�%*b�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�/%\��jX�m ޶&�hbvk~�#x}���y���>��� ӫ/��mt���������m��#�+���?}��3�L����e�eV�M�z$��P�!�A˪[	��J�/F����v�8:?�'���-M�O��~�����m��	�_��:��u���'b�'=�(J�}�֖��-�X]t$I�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�/%\��jX�m ޶&�hbvk~�#x�K"M��P�b��v݋N�����|�+��)�u��)o���r_��m����&�Ko���&�@�}7�q��J��v1a{J�h�µj�!�.M�LYq^���&�@�}7�q��J��v1a{J�h�µj�!w���{,�:g()��ikp���H���y���@�K�n�.��ɠ4�04�jfu��)o���r_��mR\�^.����c�v�J��sr�l�k]m��^~W���e�G&�A���c�v�J��sr�l�k]m��^~W���kU�����>��� ӫ/��mt���������m��#�+���?}��3�L����e�eV�M�z$��P�8>�C�?�b��v݋N������$2ܓ�A֍�a-6�Da����&�Ko���&�@�}7�q��J��v1a{J�h�µj�! ��JJ��T�zR���b��˓#���!+���}���gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�J�:�D5��h7i�a�sir&[�x�R�"�0�����&[�x�R�"�0�����s��ti�_�������C�x!�H��۽E�`E�X��WG ��l��!yZ�d/�����C�V���3��ֳ�Ե�i ӫ/��mR�MP��G�0�����:���2c�ٿzR���b�Ɔ ���Ve��˅ċ�DKY���k]m���R����{]ں1�����&.��8݄�r����6wc3�Ʋ�&.��8�,����7>���F��O���$w�ǌ߸��S�Ȍ������a�hq�М��u��9f� ��T�R��X鷴QW�w��fD���ύ���֫��XA�[���tVU�2�`M��"~6���aq��;��T����?�d���&��lΐEsE]��6�~����0.��5jDh]'\gWg��	�Z�kfc�L�C���ea�Xi��Qw�c4~Nr_�mS8<�n{R�����&�@�}7�q��J��v1a{J�h�µj�! ��JJ��T��rzj�#��v1a{J��T�p�]^�聄D&c�_�n�To�[�}�~��l*�蟾��k+Q�h'�Ȝx�5W ��̫(�3�� �f=�O�-v�*�Va�ir�4br���qP�V>t'�̗����S]�_�_��Ut�\�ą�m[���'���c�e�+���4.�*�l��=5;�a���8n
V~$�����1%��Ɇ�����5��Dao.\C�k�2v@�q	6�6]"%n��ġ��,Dd	�݌i�a�sir��=���i��?���*��4#h��z����Τ%t�8Ŕ��C������gn�=4�4�	���WdM4@��&����˶�eqm����gn�=4�4�	���WdM4@��&����˶_D⏑B[�3
�v�v-}�	mpBR9ƭ�����fx'v�ao.\C�k�Y�\��=���{&Z��gn�=4�4�	���WdM4@�肥�J�@��ey�1I0���ԏ�.fOe	�0J�ǚA���ۖ��S�<Ԣ�t9 �%�z�J��X�C������u���'b�'=�(J�}�֖��-�X]t$I�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�/%\��jX�3*��hbvk~�#x/����<�b��v݋N�����|�+��)��"L?�����G�\�4���gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�JӐ\�0�<�>��"~6���aq��.�R$���c�}���Fo|k�LbB�R���>_�C������gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�J�1�a�"O��I��jÇ+�_�n�To�[���9�P�4vE7�MW�o�>>����I���I�����OeU���(�1O,J��I0���ԏ�.fOe	� 	���R�h�Qf��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d�#P�j2E�?��˓#�������4~V��3�L����e�eV�M�z$��P�!�A˪[	��*3)�����3�L����e�eV�M�z$��P�!�A˪[	ࡦ�^��Mp�-a�D͢q��`�Lx(�i��/R#k�˟ܒ�o|k�Lb�*4��%�#o�]�ʄ�q������k&��(��Օ��qvdЧ^{�jMdGN�������V�����͹!�b
�C�x!�H��۽E�`E�X��WG ����Y꜌���k]m��Cw�Hm�̭b��v݋N������&�K�+����pP����` ��y/�����C�V���3�������D�v1a{J��d���h������	��׏�����M� �U�O��x(�i��/RŻ�&ǥ��a���F߸��S�ȌօG�j�z�2��	~����^t�zq�B&���6j�"Hs��Z�W���+�@�1!�,M�u8!n���c�v�_����J����肥�J�O@�s��M���c�v�J��sr�l�k]m��į)˰ ��E�d���8ѵ�3�L���'s{	�h�v1a{J�}D7B��#�W�/�#+*f��3�L����e�eV�M�z$��P�1:W����f�E܋0���\&<���v�߭�wۢ�L�@�U��C�|J3J����,i����׉�\�	�NiUL��˱���v��E�sr�S�
�۹�ɟ��X�G[����t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��y�]qP_���hju�{�V�Ջ~�D����zޥ�[#�P��G' �K�Y-�v�(�$�T�+V.�V
F/������Ō����<�6�Q=�Ɔ ���Ve��˅�������k�A���ۖ"'��&އ���lc�ڕ3��t�>�!�(Y��Ɔ ���Ve��˅�a-�Ʃ��_�n�To�[�}�~��l=0�� ��,����Îhbvk~�#x���D�#3��,�-��L��)܅���o[�a����c�v�J��sr�l�k]m��^~W���A3�X�N�,����Îhbvk~�#x���)kbzf	�$NT�I���I�����OeU���(;�~1��_��@Z
��#���Fi�"τ�����p��}��aq��9��,=O�nQ�rV~��s�Ṅ3
�v�v-}�	mp�r3�<q�uR�#�2��A���ۖ��1�:��o[�a����c�v�_����J����肥�JӌKa��m�8͹6���<om����J����s)x�?{���x.�KnqkH�D��3R�e��ł)w���m�±��m|J�}�֖�#7S������v�>�w�N�Er��oIIb�*���*.埲�^^V9D�4��VJΣ8#�(�>^�l��e�eV�>�3�eZ~]� ���_�hbvk~�#x�K"M��P�b��v݋N�������6��{�\�0���e�]��9�u�jsJ��U;���v�8:m��~�k0uR�#�2��A���ۖ��1�:�%�\����*\�9X����[JM�D2\1z���@qP<p��1����e��@^�11|u='�c�a����gi�Y
�,3�^�P�qjhbvk~�#x�K"M��P�b��v݋N�������6��{�\�0���e\Ԏ�=SCp���7
Kn\�H��/Sg�w��'o�un��7��hk��Y��A�m�(sH�DJ��};��*�\G�I))����A�m�(׶U���]���J6����"'��l������O05 S�s�l��_T���a�aq����.����Vc�$J�{�����~�=��K�I0���ԏ�.fOe	����4�l�>z�Vg.N������[� �I�������m��b��v݋N��������џH��zb����2�ę�u'b�'=�(lqpބ�;g�Ǣ���>���1p����@�M���g1�#�(�>^�l�'s{	�h�����-VL^օ?D^���k��^�1��dc�@c�����h��-�����s�Yls��8��GM�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2��ͮ����̩jv�^wbQh�"E&�
)H�{���8EH��q���<om����J��RQ�\Bk�	x�Hr�6w��]W�I))����A�m�(CyQ�/Ap���z��R��}D՛��W;���\�H��/Sg�w��'o�R������#���Fv�o�E�n
V~$�����-�G�h��\`�R�kA7��V ��݇!�
D�Z���䁎���w�=��u���'b�'=�(J�}�֖��-�X]t$IDW��E��q��u���'b�'=�(J�}�֖�
�c���zU�s��訌��v�8:������fI��jÇ+�_�n�To�[���9�P�4vE7�MW�o�>>����I���I�����OeU���(���fe]��_T���a�aq����i��on
V~$����4~V��3�L����e�eV�M�z$��PКą���g��j"jȩ�i��N�Na����g�6���Q,|6.o�7��g��]�J*�Rs�08�b(��R����� ӫ/��mt������q�)]Q�x��r_��mzf	�$NT�I���I�����OeU���(;�~1��_���̙�R��I���I�����OeU���(���c�Bd�����}�B�A���ۖ�k�V\�#P�j2E�?�5ߧE4�훬�pP�n���3R�e��Ӵ�"�6j��;٬sf.�r� F�3NA�׭�%*b�3R�e��Ӵ�"�6j��;٬sf.�r� F�3N�rz�f�������
��\�H��/Sg�w��'o�UX���e��o�>>����I���I�����OeU���(�*/ˮ78�I0���ԏ�.fOe	� 	���R�$D\��z���gn�=4�4�	���WdM4@��&����˶�Ka��m�8BW�R7���r_��mX�C������u���'b�'=�(J�}�֖�#7S����DW��E��q��u���'b�'=�(J�}�֖���p�5��z�X
3kZ��5ߧE4��p�-a�D͢fU�9�׏�����M�[�S�n�H�,l�����(4G��>�S���%����g���hZ�Z����pG�p�P�m��������a-6�Da��J6����"'��l������O05 S�s�l�?�D�p&��2�ę�u'b�'=�(�Y��4Q�/�5��kƸI))����A�m�(��C��AF�L�J)���wj-�s�7�����p��l� mr�m�S��^�Tj��^�G�38bS������Q���Ʈ�!�����
~��v�x�GaO�՛���|u='�c�a����g��G��n
V~$����\|u='�c�a����gi�Y
�,|�S�
���N�@E�V)�jP|B�1�`�
����"L?���N��-���'�[�s���J��sr�l�k]m��W�/�#+*f#�(�>^�l��e�eV���E㨀���:��KY׏�����MW|��6�C��(3��7�q��J������-VL�*3)����#�(�>^�l��e�eV��_�vԡ3�@�ԍ��g()��ikp���H�����V1G�׊g{Y#0����l��=5;N�����OZ�P���]��L����0�}�}�5���R�E�M09L5�>�5C'��I�Llqq0�l��Z�M*.��XEE�&����1�L�J)���wj-�s�7����4�7�K�Š��:�����<F[�z1m�I�
ZW|��6�C��(3��7�q��J������-VL�*3)����#�(�>^�l�'s{	�h�����-VL��.�I����u��ſԋ2�̙Db��E(�\�H��/Sg�w��'o�UX���e��B�`���"'��l����C1zh�v��P����=�����|$�b��G�䣌�$D\��z�
ɴ��z�4�	���WdM4@�E�RN�- \C��(3���-��w��k]m��������C��u�ڮ�C<�o|�S�
���N�@E�V)�jP|B�1��C��AF�T۳�͕������4~V#�(�>^�l��e�eV�>�3�eZ~�/t����"'��l����C1zhT
�����=�����|$�bgJXC�j�J�1���K���L���O�D mWNHN��R������3�$�������M���LQ�/8"��]ap���dE�����hpFt��Օ��qvdЧ^{�jMdGN���W���wJ���L���M?��yбC����
ɴ��z�D-'��7�q���⮦Y�m��
ɴ��z�D-'��7�q����C�E�?ݛpD�b�I0���ԏ�.fOe	�HlU�!=�՛���|u='�c�-��;��9y���n���o���*ٝ�/�K^b�;��	+MdGN���N��-���'�[�s���_����J����l��:P�&4>je`��@d:�����{~ɲ�cz���ł)w���m�±��m|f����H�ɲ�cz���ł)w���m�±��m|���~�L����:��KY׏�����Mrw�&�z<aSm�6��`O�D mWN��Ě���aT��3G�IX0F�MA���2׸�Z൝X��8�#�����c�G
�3�D Ka��p7O��*?�a�ǫcЉ�MMe9���ݱ8
l]]y�1�b�'Bee��Y"w�?��?hNp��['�O���;�M\��M���d�N-0�@��; ��=�~Y7�,����u�[��vs<��������~�T�٥��T0�"�x -�i���2���9�΀j���s��j&5��7.�ǖ��`Y�}q^J=��ڥ����Ⱦj��k�g8��p�Ǵhbvk~�#x��Og����*���[�\#���Ƹ��p��6�>/2���-��8y���#7S����p�@OM.Ir�b����g:��Ć��x��v�8:?�'���2����k����}�tM����ge���ޒ�z��6U(�<";)(F�T�M�{�|L����br ��_���cشŀ��`�z���xl%����v&5��7.�� N٣�}q^J=��ڥ����Ⱦ|����?�ٲ�F!X[�QB����.��/�EAa��G�|�+4K-��H .�/���x���-���-1?M"$�/6Lv*���[�\#���Ƹ��p��6�>��	�hSc"�HQ�n����8�E�f��5	�� ��іG��%��<�vd�̪���B)|D�$z@Q�:�T�$��$D�}���@}�%����FĪV�aa�h�Bv�z��tM]i�a@���:߀��.��~r���ř�3Y|�+4K-��4~H�<�&��x���-���-1?}3)��*��.ᬵy��f�'XĘٴŀ��`�z���xl%����v&5��7.�� N٣�}q^J=��ڥ����Ⱦ�$�!b���Q�S���a����˱f�렾���������jF�|���,��"1^LeS��`M�egUZ��U��+FF�/��i�q���"pd����v���J���_�[vc��Z�w8�PD�ˣ[Wc��|�R�]Iv4�$b��#�s�c�ؒ,�Xy
V��,���ޒ�z���t]������^�k/^���H> �([�4����,D|r9�g()��ikp���H���6Sa쎑t2�������50f
V��.ᬵy���Ÿ�`u�%m�Y$� 1���!��ۻ�F'i0�(=�oaJ�h��N�Mܲ���C�>y����iI��z�{d$,��>k�N��^��hJL��;���N6��!j�%^oe�Yy�8��gi5�k80���i"������x���-���-1?���U�._�nQ�rV��q�t7�&:�1���Z�8	J#"���&�^��v�8:?�'���.��/�V+�G����?��j:��*�O.�N��A$�P������5d���lz:@���3fEa�F��xW�U��)Qw�c4~Nr_�mS8<�n^1���^_��&7�䬬��_=���z���nF���<�W�.�P�����$��pe��k�J����֖:���g��U-�e>� {�}���my$�N���Uە������T��6\�4�@�� �-j�n
V~$e<�Ia��la��o���Z�X�#w�@S�@��NX(|W��po����Uh1���Z[;~ր|�+4K-��<�KWL�8���/�a/�o�@C@S�@��NX��D��(X����Uh1���Z[;~ր|�+4K-���l1���$�8���/��ݾ-/�uu��ڿ׏�����M��ܐ�}�|&�xVgYG?O?�v����_C|'�1p��{����~T>+��R̕q�_�D�?�JDk��q��־ŗt�K��#NWa+��إφ��<�6�@a� ��`6:���{y����i�q,?5q�p�'�� ��B@XIx�>�+X�M?��y��L��Y�5�k80���렵�!E�Y�G�˱�ߓC娤l��(Q6D���硙�t�\K7͍��|��W&":C��&*��c�fi�dL��_���/�n>�.-,��Sq'���Jy{��dN�<@Iv�H�_��Q��b�z'hۉ)��!��|"/�\�G�����dc�@c�����hX��WG ���͹�k�9��'����%n§z'�z����CU��O؏����:�xH��{as���}�pIɽ�Jz_ꛨg��U-�e�L�4�FFo*%΢Ӟe�a�f+(��SG㴊�?����q5�n��dq�8���/�"����r�S���%��Xu&�y�搲)���$:N�8.����6���zk2���dE��ċ_7�֠9�~���=���q5�n������#k�˟ܒ�o|k�Lb�5ߧE4��\�ܢ��,CZ�zk��Xs���S���m����e?�d���&���:�AS �	5 ��.�u�����t]���/�/(�[�c�eC(�55�k80���b�7��g���	0��E��("���T�\ ����Z[;~ր|�+4K-���l1���$�8���/�!,1 ��Ҟ���0�������Zm���RvT?���J��J�)����6U(�<"���[;���T�\ ��G��$[s��6U(�<";)(F�Tu�9j7Zj�ǖ��`YĮ�RUt�E��6U(�<"\����묤?���Jn�O��Ե���ʨ )o���f
+���J�)���s�����@S�@��NXD��f_%9a��}��L?�i_��ch:@aS=�?2I��� �4~H�<�&-䤔���8�j��k`�[�M�A�E�I�88s-�`8���J:��A@�r$?:K��k� ���g��^R�Y|";�!��9����3�3J��u�Ao��%U2�h=c���9�Y��v�c��Q��"��0��C��-��K�E�sI�I))����A�m�(��nb��I5�4`UV#-�[ҭ�Ă~�*o)���h�#wA֓&Zf��%j_H�ˉPM�e;�C��8y�����\�HtK���Y�q??�d���&����C1G�v��X���IQ�^.)�H[ɳv��X�b�zc0�]F:����Į��KH ��C(��~]/�f���i\�H��/Sg�w��'o¥������zP�w:Ec�[�p(	�d��;%�Ҝ���o5X�nd���/��U��{�c�Y͏���Y��)�k������o�3! �����N^���M�� ��!Z��|<;��|B�'	�?��[�bt��N&ڀM�`�TM��C�_���O؏����:.Ӊe�1��׿V�O�`���vw_���_#��1��e8�b,7��6~�$��Ly��l�7�wۤϏ�1ƍZ���t]���u%���HN}�����*�4br��\'�s�@#F���o���F�E�ϛ�~�6,�^��D����\{ف(�7�1X�iRd��D�����X���*"��Z� Ҳ́p���N��U��������U��)���Y;e�iK ����)c����_� �n=\f�5>���r���l�x��W Qw�c4~Nr_�mS8<�n{R�����&�@�}7�q��J��v1a{J��(O T'Q`���$���^��y6�T���1���0������my$�N�e�&���6X�C������u���'b�'=�(J�}�֖���
�	�v�׹��t��`�J9���_����dN�<@Iv���S
",�IC��&*��ا��=tu�w���"{�׹��t��`�J9���_����dN�<@Iv�H�_��Q��b�z'hۉ)��!��|"/�\�G�����dc�@c�����hX��WG ���*4��%�G��Hb$�wH���zf	�$NT�I���I�����OeU���(n��_l)�t���q5�n-�@�4ڧ%�fL[�j"jȩ�i��N�Na����g�6���Q,|n�@Mb���ܴ8`���r%��ɷK�� L�pMg.6�kX�C������u���'b�'=�(J�}�֖���
�	�v�׹��t��`�J9���_����KF��D1c��I���I�����OeU���(�� SU�^����q5�n-�@�4ڧ��e��t�z�X
3kZ��4br��L��_��R��n�J>|�
#�`�^{��u�oD��񔖔�ا��=tu����Rpy2:�׹��t��`�J9�������K���L���4�04�jfx(�i��/R�*�W�Ǹ���~�LM�w�r7e�e���uMV��	��y��_�V|��j(�QHL���otscC7�F��~!�ף��U��+�Xa�H(�˕�e;DOM��#g�k�����Oд�(D+R%��[\{ف(�7����n�5�����}�pIɽ�Jz_�;��|B��J�#�p�7�,��n6�o8:4�I���c�90��j��e��`���φ��<�6���n�4����]��!x�>�+X�M?��y��1�<T�b�'Be�X�;�Q��P(�R�	3i�\��׹��t˔R��}K7͍��`���-��G	�Qu��a��i��N�N-��;��M�z$��P�,�bP$���/�n>�.-,��Sq'���Jy{��dN�<@Iv���S
",�I?�.>#�����c�v�_����J�����&����˶���n�5�����}�pIɽ�Jz_�b_X�XV�b�z'hۉ)Ժ=���]�
_,vF����JVX
���$:N��@�1�˓����Uh1�b_X�XV�b�z'hۉ)��R��삅�ڭ��*���!��|�Ɛg)x�D�����X��Q��Y��-=���]	"e��0�U+�qbp@��X�H�d��JXl'�T��~��Uг�|<�9�d�L��Yu������50�����.���8y����+f�8�ï,��Sq'�@8�Qq���z�#��S���*�ey�p�?"�Ɛg)x�D�����X��L;Л���������\�.�۟���J�)��	3i�\��׹��t�M��|S�/���[�4�f,/��U��sݐ��,���$:N�t%��zxa(􆿳�e�&���6��rzj�#��v1a{J�|����$/�pX��� xh�Ɛg)x�D�����X�,?1�����C�x!�H��Tp�����J�O�=�~���=���q5�n������$D\��z���gn�=4�D-'��7�q����
�DB�%�$pX��� xh�Ɛg)x�D�����X�A%�@* ����c�v�_����J����肥�JӔ=�	o #���}�pIɽ�Jz_�E���7t�u��a��i��N�N-��;��M�z$��PЄ� *��e�/�n>�.-,��Sq'���Jy{��KF��D1c��I���I���C1zh�6���Q,|��0��x~���=���q5�n�����ŉP�HS|�4�04�jfJ�1����ݾ-/�φ��<�6��PT�!�߭y~� N�6j�"HsF�prB/^�6�\����,�ǰ�98#.�ƣ�j%�HK��Y�!}JΔ��%�Wp�B���V� ���r�hr�W�Qo�n<�!�9����v��K�@��{�T�l[�·��`�LR	9�s��;Ce,OL���9�	kٰu��b��E��'Z*)�����k!��V�_g�T���Ӫ!�J��:����N��	�Ȓ2���)5`�H��<�C�z*K��r�&U������G|M�E�����+T^���\�}�*?�a���@{2귑�U�8N#�|���P�|T�i���ϴ�k]m��v��z_QZ ���^"�R<�����á�~O�j�)6)-
����,�ǰ���9kn��회�h�#5p&P<Fs�6j�"Hsc�;���\��N�3"���ʻ���:�4��.'uy�/�8yv��U��+�XhU��`��&� �l+�8E���|�/������Z��Ջ`,9�H�W��`�z����k!�\Z��K��qb	��G�E���|�/�����y���|����4�[)�j����0��6�}�%b���2�՛�*�C�x!�H���<�n�gV��	��yvѧ�_�.�����Ry� �y&;��|B���E�t9��N�3"��h�&6B����1B�:ͫ�����6����#'@Nw���D�&�߫���hhAS̭��u4�Β��3,*��M��'��S�p��*���J�	�LÆ�c�9ʼ��$]9�(b���A
wY�����������EXs70�U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&G�'.�T���Bf����yeWq�B�my$�N���Uە��nH5��?[�O���&z���ڵ�)��$z�}�Z��b��y ��X�ıV�F3w���|���<I;}%��.0r�`�N5�Hɫm�"-G@驁��@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н��I��� g~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D���=��M\Dy����iI�]� ���_�hbvk~�#x��q��ZV��-����!�`�(i3�����_��ud8�sO�.ᬵy��=��4H��u��r��!�`�(i3�d�@���GU�lP4��/����*Q!�`�(i3�����!�`�(i3���8�2��w��kf_����d�bfĉ>99��o|k�Lb�����1%�ol��Ә�!"������.ᬵy��=��4H��u��r��!�`�(i3�d�@���G-*��jܼ�{!0g|12�mj�6 y2��R�՝� s�#���k$ �>=���#��he=��$M��DU����3
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�g��ޏ�������v��2Y�$@[�_zβrv���� �2;Β����(�ͧ+��<D'�Ɖސ���U�8Qf4�w�;���N����
?�d���&�f3s�?(쩆�w��kf�:N�B��&�}�z73$³Zj�@[�_zβrB�ek�5Wy:4����׸�Z൝���U,��X�G[����T�}ɻY~�y�����[�]9�(b���J��:�����#}�{�|VO�⅘�φ��<�6�@a� ��fFMqlgd=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^	�)��&gh^�?�K7͍��|��W&":C��&*��c�fi�d}j�����nF���<�W�.�P�H'z<�0o
zVcP����Op��V�h���w��	Ql&�Ⱦk���4br��$��x�-n��>�my$�N��]流�>���ݤ�E��p�$g0�9Ǐw��	Ql��gmJ/��%Q�[�J��]�U��97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��1�m+�D8�̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н�QV�=��̟�1��M���R��ӟ-���J��RQH�RtV�^�'��o��̟�1�C�|J3J����#�=3!�`�(i31���~!�`�(i3�YN
��)e�'DV���b�z'hۉ)��d�7�q�!�`�(i3�5ߧE4��!�`�(i3^()��>��VTҝD!uǴc�1�RG�p�P�m������� h�ҩΟB�'��a�S���%�������VTҝD!u6 y2��R�՝� s�#���k$ �B�'��a�S���%��3|v��Eb�z'hۉ)��d�7�q�!�`�(i3�5ߧE4��9�d�L���`�����G��Hb��a-6�DaM-��&ほ�dE��Į�Ц���Օ��qvdЧ^{�jMdGN���M��ZLh-S���%��V�c��ݘ��o���F�a�D��<?Y��Yf�>je`��@d:�����{~�
\za$Ad�
��9���>f5�� b�z'hۉ)��R���p�-a�D͢q��`�Lx(�i��/R�K:+>&aD�4���t]��� z�P��n
V~$����<;@{�t���=�g��M���R��ӟ-���J��RQ�%�z�J��
\za$Ad�*8Җ�N"�g~:�âq�t�d4��W+���xȀ��D�[b%Ɨ�g����Ǵ=q@L����,I&6{~��e��0�U+�qbp@�3t���=�4�04�jfrw�&�z<aF�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��#}�{��Jw��3��.�g3Zv���� )�W/πs����N�KRK���DV4�ސ���E��'Z*)�?�R��n��h
:h����t�h��W+��W��4br����'�QV[1��<[�(yJ+���n���E�i��4br��yO{��`�
n��>�my$�N���Uە��
\za$Ad�*8Җ�N���C�3rEe��0�U+�qbp@��.�g3ZB�ek�5W� hew����~͏��ޡ�m���Y�$�����"?��A$�P������5d��n4s1��7�癆cgQw�c4~Nr_�mS8<�nt�{#	�x��Z�8	J#{�N<'��I�y��!�P>�h��@�19TH��6�!˓C���I�Au����V�hdWk졾]wL�CK)�yy ={�%�싂�nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r���Zj���
�4br���qP�V>t'�̗������^ā�Ӱ�|��v��P/0G�D����M��p�#���Fi�"τ��X��WG ��#��۲�,�y����iI�(�%d�#Tzhbvk~�#x��	���1tSjv�!�`�(i3�͵�p�w���>�$�݋\����>�������Ra])n#:�����{~��萬��]�p� �!�`�(i3��Ě�����}Dq�f���Ě�����9������n)5,�O�޳!?�R��n}�����H��B� �b��!�`�(i3���$��@ɆJӱ�z���=�r�l��=5;�a���81tSjv�!�`�(i3�}D՛��4��"�c]p�5�	Y�F,p>)!�`�(i3�šB)���4�zB��ɆJӱ�z^օ?D^��!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��rw�&�z<ad,��B����,l����0��d�����4br���G��9B �Z����pG�p�P>M_���Ut�\���ii���H�w���^�×�umn�q��J�)4���δ��;zQ뙥�X��#�^�����K���/�ciJ�h�5,Wlr�r%)cA�*�gl�&x�K:+>�}D՛����3S�s�A[��E};l�-�����ɒ��n
V~$Mr��p�ԍ�S��4$:��{K·f;[����"L?���1�����Ǹ���)/�~�T���]'�^�����P�HS|�4�04�jfB�R���>_�u��XC���}D՛ؤ!����'��M��2�B���l���_wyt��:����
�K:+>�}D՛ؤ!����'��M��2�B���l���_wyt�J��2���$D\��z���g:%���5�>�k�FTuءL�\���:��KY�[b%Ɨ�2b���J����w_���!�b['٥��gV�J�1���K���L���O�D mWNHN��R������3�$�������M���LQ�/8n
V~$� ����%��>M����?"3�m�����h�Ѽ�o������S����4br���qP�V>t'�̗������^ā�Ӱn
V~$O���6�[�Sx��ۍ���#8��c�Z�~��a�z6��}D՛؊,H0���-��M��2�B���l�2��Fm�ӫz�Ζ�XƤ5_���M���R��ӟ-��濫�L�ፎa-6�Da�N�]�B���vE�fc��57'٥��gV�x(�i��/RC�=�+c�w��9��4���;��%YX����A.�%A��C(Q6D���硙�t�\�N�]�B���vE���GFOg�S�<�c���6�N�T�\ ���:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vx�m|���{���{�=0�E�ϛ�~�6�!˓C���I�Au������h����N�]�B���vE���GFOg�S�<�cث��c�3e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc7���8��ƶ��^���R�-$M�4�	��r�j��V�������1��\�p�������L�1
H�3v����f����T��� �S��t�P�4�H��5��<�>��u o���*�|lCY�o���KU�M*��a�b��T�Q5
TZI.(sn��.u}-`e¢Qw�T���wP�|!�`�(i3!�`�(i3^��	pM��^]W3��Xi�H�=�d�V���G�8e[u�;0�ht��p���b}
�QL�����:&�ĶDT�\���wt�퇼y��砒���
�r-����\��/��WcprG�&[���� 1�Hl��5�9߫�%9!�$i�� �4�D���@|�����Q��I3
Α�^�*?�j�F��?�[4ǿn	N� ��{9�%��p[��������Z��n�G~�,��8�1ޞ��&e[u�;0�2����k�Ps_*�GqW�w��fD�]�K�]o�2�u]B>���ć+叔��r�b,�
Pн�cD&���ʰ�E;Eh	��Lx�A�B����#8����쨷	�W��<+�Jg����n1�;/�6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3����]dF!�O+�|/������Lx�A�B��8�nb �z�g��U-�e>� {�}���my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&rG��Hb� h�ҩ��T����ML_��f� 1D���M6�W�.s��錛�%`RD§B ����z� 'J��@�D�5�>U�m�j*��{�%L_��f�����,���b�������`y����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��mךBo�NgC��	��KC���?����P 'J��@�D�5�>U�m�j*��{�%L_��f�����,��9VP�=1�<E˞��DV��	��y�i��3�%�Z�Xp�`�<�..�4���ho7L��2�"�G�p�Pڹ��/^�w?�d���&�N-Y&yo�q��=m緒X�X�pF�{_8�Y��=�}�VݨyY��0Kqɔ9Q<ϯ���쨷	
P���ɒ�!�6UVo�˱&A3l|����"�`Ec'�\Y-φ��<�6�@a� ��fFMqlg8����z�:Fa�7�����~�Lk݁ 1���tw�i��scX{�X!,���{���#�0�zG�������&G���y��lDtD3�:D���*(H=�ƍ2���l��^{T~H���^a�nu4Bޗ��jw�	���ݚ�Н���fCI��8��GM��-����!�`�(i3S�#p�ۥ�Y�m#� �,W�+�dr���ͮ� л��5ߧE4��<�6�Q=���F��O�C#/<���q��ܐ�}Ĕ�ttvfs;����^FF�Q�f���S�$7������φ��<�6�@a� ��fFMqlg8����z�:Fa�7���W"�P�K¨}�n/�J� &�0D��R���Xc�Qw�c4~Nr_�mS8<�n�ݚ�Н�T��a⨯�d��+���{_8�Y��=�}�Vݨ��}Dq�f���b��~�F�KD�Vr[/}>5��0�B� �b�в��y��lD��KJP#�d��-��!fM�N$r4������8!��?V�&�2���)x�?{���x.�Knqt�dĳ�ߗ�ݚ�Н�E]�tM1-����3R�� ,��rQ͒������ݚ�Н�烉s)�v�bP�63Z�t��Qѳ$G��A0ok��烉s)�v��IX0F�ML��M����4�	���P���/��.�g3ZE��g�Hby���=)�Vk����/x �i�{��R�S��>j���T�}ɻY~�y�����[�]9�(b���%�fE�D�8��w�=�-�R3х���W���Bm�����y�3t�ʨ�u���C\��~g��tcb�A���t�T��?E-h��`f���s����a���'���_�)�fo��&�[zL͊�q���\��;�,���+�^n=\f�5>����Db^<�..�4���x�H@�[\���F�`yx�>�+X�M?��y�!�`�(i3Sm�f�e��N�eM�#��}Dq�f���NƥNoz��KUq� ���F;p�	�	�����e��0�U+�qbp@�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r���'��o�u:��_x���O����]�!��	Ǹ�y85��8��,	iL�*dgN;ۍ����$9���Z��o�^��D���:5A��p��(1l�jG���Z��o�h�G KH�F;p�	%Ɏ�Bi!�`�(i3�ݚ�Н�-��)'���N�R���Va�irl�
@\�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н�ҷ��.Gɔ9Q<ϯ״$(�>g�!�`�(i3/w1z��ӊ+�`R��ӯ�2�`<!�`�(i3�d������)���܇�b~*��s�OY '��M���R��ӟ-���J��RQH�RtV�^�� л�����P%��v��!�`�(i3uD�*'D��?�$���}Dq�f��	��x��ݚ�Н�ҷ��.Gɔ9Q<ϯ���쨷	
P���ɒ��[�a�������������W�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j �_�ȇLШ��+���Al+�H)Z<��n$7������φ��<�6�@a� ��fFMqlg8����z�:Fa�7���W"�P�K¨}�n/�J� &�0D��R���Xc�Qw�c4~Nr_�mS8<�n�ݚ�Н�T��a⨯�d��+���{_8�Y��=�}�Vݨ��}Dq�f���b��~�F�KD�Vr[/}>5��0�B� �b�в��y��lD��KJP#�d��-��!fM�N$r4�/	<ԣᲹ!�`�(i3���w�ze���M���X����Ľ���:/��N�g()��ikp���H���Zg(b�d�w���	�e��D۾���!�`�(i3���w�ze�4br������Ľ����Չxv��Օ��qvdЧ^{�j��@�
h����Z>ؼ��XyH�RtV�^�G��^���J��sr�lv{��lw	!ݞX�����}Dq�f���Qѳ$G��A0ok��0��l!���O�D mWN��Qѳ$G�φ��<�6��}�6�nq�4�	��"|�1�2[u;��|B��loXB�R�S��>jȅ�zn8J�6g�#��%m�7s�B7JQ��H{���W�.��A$�P������5d��n4s1�U��B��-";o!��g��Y#&����"sS<�0�zG�������&G�N��W��pp�N1U�)P<�ܓ�Y�������b@����7)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G��+p��qR���Csht��p��^�#g���
ۼ����g
aC��e�ݚ�Н�ʬw�S���<v�cn@�q���uҽfĉ>99��o|k�Lb��Nh�=f[u>a|��X��WG ���p����[{�o\s���x(�i��/R}�	76�&�� Ӗ�t$�)�vx�؊ګ�$��t���������� �8K�v�~^���H> �B��p�b�\��K{h�I@�?.��N[jX�.K��o�5�[՚1Dq��P�<
����}�Fe��1��dJ�5!�_H^��Ƨ�0͜��!?@K�F~�����/����ϣǖ��`Y�Hw��pZ��T)��>e��k�J��^F�=/p�i����T��T�^���h�.k�mb�&��ƭ�����Ǯ;����@{b62�tstF�!��c�/�g|��0.����;qX�qp�c� �����=c�!{p85v{��lw	w�����!�s�ˑ����Oh~�o��_�Rv�䩲$��V���,�wOC� $�0�n=\f�5>�V�/e�,�G�6iX�P=��HF�9�Qw�c4~Nr_�mS8<�nC#/<���q[�л���7Cw�Hm��K7͍��|��W&":C#/<���q*qA����6\�4�@�� �-j�1tSjv��*TH�SO=�O�-v�*_�mS8<�nC#/<���q?V��j�c�'�QDn4��F�(=C#/<���q$f��_Ub�}Q�sd��fINY�"}Q�sd��#W��r�S�C��-�!� �Qܤ�6�W%�*��Rl���sp���md�g<I����2�"�G�p�P�(��Iw?�d���&���^��[� <{>w�\퍜��Y��>1Y�V��	��y���x.0��+�Lw��riQ��[9-|���vG�E�xc|�'�6��Ĥ���M���R��ӟ-�F���ˏ��Z���G��^��k݁ 1���tw�i��j}��wF�36�o8:4�I���c�90B3v�A��ʃK�,��`U��B��-����A�;�����\��]8��	�����;c�~5��IM�Ex�>�+X�M?��y�!�`�(i3��Vvq�#QSU:�����|e"@20߀�5����.��	�����e��0�U+�qbp@�<�6�Q=*qA����6\�4�@�� �-j�1tSjv��� л�e<�Ia��la��o���H�RtV�^��Q�Y�t��ܜ�[��H+�����'�,�Ϫ�!�`�(i3��z�������}�Fe��1�:��g�XW�� л��5ߧE4��<�6�Q=���F��O�C#/<���q��ܐ�}ī��K��M�ZP�����Fz��Ԥ���엝�����L}�]���4x;΂��m9Ϲ@��2�{��jo�W�ք�w�xW���s"�J���_OB,8��R��TR���L�BZ�?=:�A@�G�PY��Β����t�T��?E-h��`f���s�c�n��X�`���φ��<�6���iE,�p@٢�ԡ�p5��IM�Ex�>�+X�M?��y�!�`�(i3�>8u]�ZL�q9+t�}ȓM�Me���`6X���dc�@c�����h��-����<�6�Q=y�}�6f&rG��Hb��Wv
*Tȍry��	�� л��`}��vv㪤�vF}���V6�pz����ʳX��9������yi�@��������zȜ"��X� 2<�6�Q=c.F���Z �W�VL��׬��P�|T���nT����
y���^��D��G��q"Y��;����rx�pj�d!�`�(i3��ǻ��nL���B��6�<������NM����� л��5ߧE4��<�6�Q=���F��O�C#/<���q��ܐ�}�2oY��.��Qѳ$G�;��|B�dj4��h��zɾϞ�E�md�'1DK�����QQ����"?��A$�P������5d�y7�����iI9�o«IX0F�MR�c4!`{ਃ�6���po守�ubs��2[�a��o���H�RtV�^d�'1DK`�I��Wn��>�my$�N��o�/���;�� л�������k��O?����'DV���b�z'hۉ)��d�7�q��^{T~H���^a�nu4Bޗ��jw�	��ȓM�Me����KJP#�'����u��r��;�E���Ή~��?�kv��.V��:���������f+v�k�@1����2���'����u��r��<�6�Q=Q١Ӿ�$�̟�1[Hfƥ�QY�j�`M����M׮� л��5ߧE4��!�`�(i3���?��$,K�9+�/���p���&Cd�c#��N2D���a{�l�
@\ٟQ��ǺΕR��ӟ-�$m!ݷ�\�H��/Sg�w��'o�*0��}�+21tSjv����y��lDtD3�:D�����-ќv�Y_�R��D厺��+���l�K�>�������I��Yq���k$ �� л�������k��O?����'DV���b�z'hۉ)��d�7�q�<�6�Q=���F��O�ȓM�Me��&[�x�R�"�,bxqX����F��O�c�ˆ�A��߸��S�Ȍʞ3���h��[���x�����$,K�9+�/���p��\��be�����E8R�c4!`���U�._����P�|T�ݩ^�H(�BM�ܤm|��B�=9ODR�c4!`�d>�c�n��N.�6����c�+��!�`�(i3!�`�(i39�O��F���{S'��Sm�f�e3�� L+��M�{�|Lɋ���)���O?������T���b�Bϱ�h�5,Wlr�r%)cA�-��h�m ӫ/��m��?�4D+%�����
`���zՠ�����Z>��~��l�7��;s��!�`�(i3��7I��٩h\K�5~�!J��/٣��q8h��^�Q[M��M�ŗ\�'	�?��[��ZM������v�E���a�e56<�R�<<�U���+�J���q���U�C#/<���qHe�-�c���{L,8���Ο]_Z鎬����A��:6])��[��x+%��6��8�ʪ%��1�d�٣��>����C�V�ط�aFmғO�4}�G���n`5�fK�\w��0]����v�E���a�e56<�nX�8jg2}-}٘q���U�C#/<���qHe�-�c��3E M0�F�T��BZ鎬����A��:6])��[��x+%v�-���w:���z�Ji��d�٣��c�A�L'Qī�*pY�M�l��S�J*�Rs�08�b(������l__��E� )�&��"X��[��Q[R�7�z�C�f���Y��¤լq��/�NI����&�ߝ��e�4�+/r��bQK��Ņĕ|G���8����z�<;0V5���ܺ���0�c�S�u. �����n_��Ď��J鎉�����3[�u8�Z��}	��ۼ��*0e�El����ؑ���6�M���ʄ<�6�Q=*��^�"~H�𕎭own�~]�g����A��`-���y��lD�Vf�`H�jRj�q�wxo�~]�g���[��}��#J*�Rs�08�b(������l__���#���,Wc��Iu�RV��,(�
4��c��^�
E����d���m l�o�&�C�/�s�f�I�<6��$)K!�`�(i3-��iW��
�!�N�".Œ<�6�Q=҃���),1��m��x!�`�(i3-:��M��&�A���ۖ$����nQ�rV>Vͭl!�`�(i3w�
��Ǽ�aS�>
!�`�(i3�M����v�v��8<e�� л�?�ᒹ�G�!�`�(i3!�`�(i3���BjJ�l��!G���� л���5@~Ju*k`Ë��!�`�(i3�F�7��Y�
�cc�V��ݚ�Н��D���R]���R�!�`�(i3r� ��i�(���B����_T���a�aq��G�n���t�;���N҅�����<�6�Q=�V��(��sW��|E�q��w\F��G8T�w�nf�?ǉ�=��K_%1��x��~iM5/�S3 <�X;p`�M���ʄ<�6�Q= ��ߕ!�`�(i3!�`�(i3�G8T�w�n�ݚ�Н���u*�C@�g�o�3�����t��˳3[�u8��X�4���	A�/ї:S��I����yP2Ni�~�ݚ�Н��;�k�f�!�`�(i3t�%�Z?��<�ry^�}];�SS�jX�p!C+Tl�������l6�O��(���*-�¾L��8�$��`�� ��M�#f�?ǉ�=���E?��c����L�{��%ў׫>V��2G����j����PJU���˶��-�-��3E M0���M��s,�<�6�Q=E�%�� �-��v�-���w:7�sq֜�H�� л��G���X;p`��8
�[����L@]HSϻ���j��M�Mb�:u�!����3���3E M0�~�O��������y��lD�L��R4��&8�,�R�Ø���Ko��1�� л���oww��X;p`��5�j�))��<���՚Z�,w�D��ng�.��R:k�ڛԀlY�{:fh�3�w�	�|�s_�oAA�Wc��z�Kl�u "���
w�u�f���!�`�(i3<�6�Q=�D-'��7�USe8ӭq��P�<
0��l!����B�r��B�t�x[��,U�ߑrf�����4R�&���K�V��Y�uYu����/�e��<��(���B����_T���a�aq��G�n���t�;���N�`���EF�&'��Y_�C#/<���q�>8u]�ZL�w,���<ҫ�5���u�fJxL������@ջKf�P}�)ܙ[�@��\�F�Y4�,�<�W.?��!���k��iE,�p���6��]'\gWg��	�Z�kfc69�#��r���+�^n=\f�5>�.F<!W���t�㮫��po守�ubs��2[�a��o���H�RtV�^�s�eШ,iS���l�
���|e",�u�S��d��JXl'�T��~��Uг�|<!�`�(i3���9��ۥ`�M?��y�!�`�(i3�s�eШ,
feq����ǒÍ����d��]�Q��f�_��BvGޣkQ�A���ۖ$����nQ�rV�}!�@�?0��,H/����\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh$�)�vx.F<!W��p�k��|-��N�^q�Gf�q�	��cO?E���YPx?`�D����$6�@�ʷ	���M��p�#���F�Q���*�(S�ȼ�{���ў�L��jVѭ@!�`�(i3m�͎�=Ni�D%�<Ȝ���,�ǰ	M,��rER��k��E�(㷾���E.t�