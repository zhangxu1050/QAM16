��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag����pH��q^��+o�7\F���r����&$9g8�M>PFWD#�z":���ӳ��_�x�$t�`a\�R�F*}Ø���K�ZF��W��`k�ZV"���:��#tC���,?a��Q\�_qť��[�޿-ǋ 4�iҡ ��d�n}K-J��K��z������3�z�ω�C�I���7�	��.'���F72��{L�8br�.�/�d�������4�;y��v-.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c, '�yN�210�|��1�@��cOL`¸[
ϊdl�E���2Ee�Y�R2
�I.��	���
��i�S��/��5[��̔��o�^���~�CxT�Z4Y3>���~�)A�t�ە�.U��B�?���@���%U`g!�� f2�}�ꦃ1d��:��{�}����V�m��ˁ��l�t�|Hƿ+����س���c�B;����̢��əMO�<V�9u	�1ծ���j���v���Xt��+Ǌ���zϻ�z������Ӻq�|��U�h�r���/E�CԵ�_�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Z鎬����@�Q�2�s�JFAa�ߖ�g��o�4��?����DNZ�j׫���?_W�\I��ఽ��`g�5��!08�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"�~�#�B7�aC�h�>�N{a�9Ow�Y��k��ı��*���q{?d']l�+�ʛj�I[ b�����,\ަ�It��;���:d#���>잣����i��E����F�'n�^0o�0��wU�g��Q������4��k�y'��a��u*K6H �i7�sp>g�?o�x^[��
Bq0�[X�b\g�##qYw�J��g�U�/Ax��R�>(�I��P�O���������G����<E�ªY0�Б����!�`�(i3"�,�>E��4];ˍH�,t����t�i�lK�軧:pPFy���U��!�`�(i3�E����F���8�TP���{��XT}u��Q��eF� $���v�]wɭ�7��r�=!�`�(i3N�By3��<�]�!����M[��Ǣ)�k�4�U!�`�(i3�����5	���]����,�JL����?D�8��R�����!�`�(i3�����5	���]���>����CΌh��eZ!�`�(i3Y%T��BPe.��xu	�>��l%i�-�5`z��s�Ƀ�?PA�':E����j���0z�cUL�I��6���T�\ ��:E��]��8S�n�(�a�x�f7﹏N�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�����5	���]���>����CηxmQ,ۘS!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FH=Y��@�E����F7G#+��\w��0]�o�t��F�e{iʖ.	��A���TD��ό���.Ӂ��̰�!i�q8�2t�ݡ��1����(�
t��Y�{'%s2�ew�a(􆿳����^���(R\֎u�,��7-�)�V�3j@IE�U��>��l%i�-�jo�'q�!�`�(i3�E����F7G#+��\w��0]EOJ�uxm�j��O" w�"�,�>E����-��%M�rs�i��;m��"xd#���>��CyW�f�tR�wX��q�\E��0�Y$�J��;!�`�(i3��(�
t��Y�{'%s^;$v�P��<�4�����6��	���`y���+Ќn'I�+��x�v/cs�x�f7﹏�����
L'���XwI<��f�E�#D�����Ә�N^tӱ1R�m��+�<4��ˌ�ň��h��<�..�4��B�C &*�����R$b-iu�`���`�+N��1]�O�>P�2-i_��2�e���]/�fm��+�<4��ˌ�ň��h��<�..�4��B�C &*�%�}< VW�F��-ֿLE-L [�/��$ʖT!�`�(i3�d�٣��4�5_�o0b!��u፨"���Q�U!�`�(i3���+�J���q���U��@����gG�5�3��PB����A�E����FZ鎬������_�,��LE-L [��ak$5��f%%e�d�٣���N N�S���c��:KYЙMǿI?RR6��-z�n`5�fK�\w��0]b!��u�D��u�(n��������+�J���q���U��@����gG�_�H���	;	�J����-���Z鎬������_�,�;�7���c�5��(�Vާ���5��d�٣���N N�S��+\�g���8^�Xe�!�`�(i3�n`5�fK���ġC��װ�:�iԟ��=��.wd���/�t-gx��P�\�<��R=p���W�.�Ӂv�u�o�\�rG�,r�.!�`�(i3jݭ�F���X+�f�f�!�O��1���Sns&���)�δ��}�\���;�YǯXan��W��u�L5ӥ���98�
x�?���~46��E����FkѶ���� �G��:�lL��:�iԟ��=��.�.��SW+d�.�Ӂv{�G��ͫ������:[�F��#������+�J���V�L�X븊.�Ӂv{�G��ͫ������:[ۚܖ��`��AW˟����V�����lJ��I��p��mK�������T�-07���wұo�35DEio;`&x�jop8��Ǥ�X��1�\����iW5j��ts���k�%�(�[U<o^.K�}gm?2�I��6�]���~߈�&{�ո�UfG���$��Xo��� ���Lkߦ^Cg��)JHn��z�Tp(��v��9gP�U,��!:�ib|� %ݓ��E�v���bQXX��bF�Z鎬������_�,��i�p��+˞j��&����Q]� _ό���.�}�
�?�#l'U:�g[��爤��d�٣���N N�S��E ���� ��M�#зq8�Ј'���Xw���,DFmғO�4}��oww��n`5�fK�\w��0]b!��u��8
�[�����.���5��]�!����w�Հ��a�e56<�nX�8jg2}-}٘q���U��@����gG�.�>��͙F��6�7s�9���o��S8��<�J�QM�h���J	�J�y��*?(�QNȮ����`y����@����gG|�w��DK����$���7s�9���oC�M��N��.W���ۗ36��T�%Gvx��Or�[�]�!��RY���ت4�6@|�~��\��o3� �~x�
!O:0����-yMc|��ޯ��%װ$��_�)v�_d|��{�R�$�V�<�xwu�P��j
��rR>ݒ��lFh�]�#��mIZ�q�cݵ�Ǡ��R�Íķ"�=7�7K�Pe���b�׾ŞWsuzS�n�(�aDF�������l#-����K8�����JC�� W��$����>&S�XQ������;2��h��`�!}����U�|/r�����qȌ�*���-���*�ߑ����Њf��S8�YX�s�O����&{�6�LbE���jVѭ@!�`�(i3!�`�(i3�N��W���tRs�:�I����hoDy�����O̗A��{�W��L��x!��G-�Xy|�W�����6�BQ���4���%?K%����=ZXR&ad��_��.)<��O����&{�6�LbE���jVѭ@!�`�(i3!�`�(i3�%ؙ,{F�2������x�f7﹏s��m�Eq��`<��*�[�g���zz��c� ��c�t����Ы���y���!��R-���}o��Xy|�W��t���˵]߱��qC�G����]'\gWg��	�Z�kfcM��fZ� ��b�FP&�J�'Ƕ.�I�[�� '���Xw�j�7��[|��;�W�x+Q�*M	Ƶ�a(􆿳��_�"ۆ�}��HN�=m
��l��"����/����(��a����إ�n4s1�U��B��-|k������������r$ɓǉ�.y�U=������&G�������8����� ,�u+c��q9+t�}x��7��S�n�(�a_1�f���k���������|e"�J�'Ƕ.N����;K V����(K7͍��|��W&":x��7�֕iK�D�b=��p�:�k���������|e"��)�δ��Iћ<���I����~u/��kOT(@X~�H:������宦%��s��u"���ܹ߆�p�h��d��JXl'�T��~��Uг�|<�d�tu����=ZXR΅;&�_��9�+��N8�����JC�� W��}Dq�f�g�G��0RR6��-z׾ŞWsuzS�n�(�a�e>%�����J�'Ƕ.N����;K V����(�À���S�>���X��@5���sܑ��y���8���/�YZ*��zʐ����WՁ��̰�!�Xy|�W�(�[�*�ۢ	:j���k¶lW�x��7��PB����A!�`�(i3��X�zl�rx��E�x��7�� �����2�w����6��j��8Tʈ�Ym�����xb}�	76�&��A0ok����)�δ��+�qy�t��{�!��À���S�>���X��@5���s}v���۹��׹������-�mic�y���6G5_eOu�X#*ݔ)P<�ܓ�YV�=���i4����]઱<���E)��Iiz!�u]�MP��(R\֎u�D��u�(n�f��G� ��M�#�h��N�M�����K�H;�.��1���,:&�����qȌ�*���-���wl53�e�%^oe�YXgJ,�|dq00����M�{�|L�8�YX�s�O����&{�6�LbE�렾����k���*�Q+jq����M~�̀RR�7h�,b0V�u�Q�������Zn��޳Q�4�gX����cl�"��Z�Z�F{/����MB�8"FeIN"�-���0�i.�9�e�MW��Rj�q�wxo�~]�g���a\;V@|Xh�hk�g�l�&�͸�!=.�
kZ)� [��v���Q:�7-mł(��gR� �ұf�?ǉ�=#B��F�!�`�(i3!�`�(i3��*�{6�����&!��ȁ��;�<n�f}�T�NHX��+���;���5��K��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3w4�4a0E5' �c҃���),1��m��x!�`�(i3�(�;��NPf�?ǉ�=m3�țZ��_�`I� B�!�`�(i3�<��N�Lf�?ǉ�=?�ᒹ�G�!�`�(i3!�`�(i3���BjJ�l��!G��,3�/�r^w��'�k�f!�`�(i3XO����0d#���>���6%�as���eZ�c]��E���!�`�(i3Q)��Zl���w���4Wt#�X�S�n6�P�CQ��Bރ;�{��C�{����K�7��(�mWƒFR�6�!��&t�ND�������K�7��(�mWƒ
 ��4���>�*�!�`�(i3���K�7���]�i�hv�)?`��BH2l}�{rcKE#���.�)�p�ҀL���G���ȍry��	X+&wG��	-�����8�%�b�-�#G�<�ry^�;7hZWT�-��$ϙRl�bu�	?�cx��s�٩��!�`�(i3���*[UxG�2��}����a#�f�����JQ	�c�kj� #��� !�`�(i3��%ў׫�o��LD�x������	A�/ї:S��I���fÓ���(�6k�4d��^�v���/ӳx��R:k�ڛgf�mk�*��^�"~H�҂��hWj���H�D���dݮ%*?�k�V�?�҄���>�8�$��`���	(��7�f�?ǉ�=�G���X;p`��8
�[����L@]HS��e�MW��T��b9���ey�E�����$���f�?ǉ�=��oww��X;p`��5�j�))��<���P8C6k��\��ކ��[����