��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htdʮz_�0�`��@�[D˂8��k�ľF�n�Ԥ��r�τ�u�&&����\l&�$������<H�����}�ƌRS>�(B-~�� ��ڣ�9#M��c��&��C:��p�����>�.��`��*��(���P�^Ս�.���,�-����8'bɛh��7�8_s�o��7]�d�7�#//��l����_���:D��u�ϩ��x5�qܦ�j����h��L�&-̥_7ż��_�Xy��}S\���<���u	��p7� 	a='�����i��Cr�=�mP�p�9�룭'��C�WZ�4�A��1[o{�RϾ��!�8��������@��~OU!�U���,��a�n��4�H�	�>��T�a�P?Z�w�}}�;�Y$�0��X���I~�A�wn�`]XΆ0�z���a3���w�e�m���^4�'�RIQ���'-W�d��RޏvG����<ޚ_�y�Do�(�hf���KYf�H�6�u]�щP��5jG�Q�^I�-�ø!�v��;Aܦʳo��ą]T�S���G�:v��V�\1�֖p����p+�	�^=�1*�洘��\�.���X��m�Z�
�$d0,�ֶ��+R�"�W�9�����U=��u*W$�
1�Q��b�4"��p~񊥇�����s ��x,�<�HaC�̾wG;��N\F!�i��T�T=�r��!��t��7|4ay?m�Lң�T_\ɝ��!M(�Y�u��N�*���1�ѡE�/�H��u�{5�6���4Z���E�0N:p�k��e�Kk�����ׅ����)�}>g�Y	�����.��@��VV���j#�O��d/@xp"�S��N8x���U-nR@.��&��݃=��U& ŗ��j�h���c�d��osK�{a�0�[3v�3$�\w�U�!C/��,��8���%iQ�*a�bB���|�����U�,!�#J��!���̓m�D����6e>����c27��`�H��d�tu�=wZ��J�����x��D@�}�R�_�R3�ӀГ��]x��wt6rg�5j�4��X�M����R��v�%F0ťƑ��o��2 ������>^em�������omi7{$��m_�2��8q�3W���N16�k�k���~#�gfyٶ�}�?#�A���xF��̐vži�B���1\�`��[�v�� /kJl=Jy�� }b��aA6D��x��.�i]^%�&�%�M�����e������-��I/�G��}}�]B���31@`;=Ѓ72�A��� ����&��K����>���͕�U�����f�����BQ���M�U�o����Q���~�Uj}��fTe�F?�w��9ލ@����@�qN��J�{���\p��< }�ys�,�3�&�$������ �Φ��(��V����Dp�ȱ�S�Sl��i"�S���&�e�L�~KG����.Ҍ��D����IJi,���%�rc�5�v|s��KY ��p.%Ώ��W�B�.�`�Re9��\����"��6?M\ ?��&��֒/�R������0�PU+�P/��_�:���rx�59rq�^����=9�3PvԽ�GA�^<U���a��4I�Hm`�뒉E�h5�dE���5���ҋ���5���؝��9}b��+�EA��#&"?�J��P5�)ڂh�Y'<����4�/n}g�6V�OmYD+���(��@Щ�*��V%%ҩ����i�s�G.������QK<p���.��UU򱖒�Y�_�~|�$�/q�2�˧� )�1���R�^ٖ��`��.�A� >�5�I��Dn��kJd�+��p�����7��%Mi�~k����Ge�]V�jv�^B-D�e�ܧُ<Ͷ�޴6.P�=K��=}��?��D7�/�����UÂ莟bӧ����k��+K���v:/�c|��&x�dp�wG
<�0�8��:J��Z��+4�L�A�����8K#�VƪV.���z{�� @��ۧ���`�%��2xNT0s^� ��~���S3
�r��]�5�+�F�D��d��&O7[_D�ތ
"�z�^�ɷE+	�*ťX��@X���g�"q�\�*�0�r8F��d;6i$W*���NB攏��63��8�ꜗ����[�cˎj��q�N�����5I
���r�/��-}n���-k�p0MPPSn�8�ZH#V��P�'��~M��姺�,��I��p�疹k��6���e6Z>�j4�� ��� z�]��%��k��������خ
}S�����y�+-]] �J�$�6�KiU�y���^�V����~N4TE�͂�6������N���RO�S��c��f���yj0+
�C�b�J�9~���1�U�r�}ۖ�}��ĥ�i?�ҧ�h�H#"�m�������X2@�2�1a�L�6��G�U��E�W�cQF̋�}�lf�U��i.Wxe�ˌGX��&]ɞ@��I�KRֺ�DG<�jC�wHr�1 2Z񶟇˴�w��l�/
4��h�摯�eӪf��~Uq���D�M�挃=����$�0M�r}X����;�\���Q�����Ǹ�!!�"�,�0�o�|n��_g�Z�P}����=U���ВJ�����f����̸҅�<g^K��TQ*A��la��@.�8O�	�GU���a��2HK�P��i�2�%��K�b)	�́�	����'�:j��ʎD0�#З�m[��`>&Vw$�\&Z_S�h�30�0,����}d"!��\�v{L�^^)�G4;%
�6-���]fVD�}�Ʈ}��0朎�x)<�-+�k����e&�٢�V��lQQ��j�m��G�}tJ��!<�톢y��p"N�6}	��Ī� \�L��@}���kGF�E�t*�s��"�"p��\}QˎZ���X�Mi��b���K�>�S3-���+8�*��i��O<�CP�^�y��Z� E8�ԩ�P�%qh��c�z��Ѽ�haw9�����<it�h���P���r�9��)P9���#5��4KtS~��N�6dP>D~��C�B��V��/�\�g�V�mn��ͷ���˙��8��x����A[��P ������,��#�Xެ���ja��q2m+�b���־@�	�%,�:���G\9�AFOC����<I��F+|��l��z���A&�����P3WV���@�Sv��g�o����b���y}J!$LO�G�u9���[o\���Cit����xiwnT��(pL�