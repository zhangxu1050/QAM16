��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR��OMQ�bs	�.�z,yN<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR��OMQ�bs	�.�z,yN<��;��� B]�pE���	x]̃Dj#^Da����M�Ov��12È�pT�7y��z����)�,�˛D��w���旴4�����:��@���b���$[G��m$�;�`��v��p�㈍x���t�켻�S���c,31�-elwB(�93;2���Zߧl4���0�?�1~�x�c�>j����d��S�W�>��Q�d����t�mR��:�����-��3���7�Jk")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc/?�s�m/C�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEA�i�+���Y�y��
r�)�Y¹w����i��T!R����.�D���J7"�~�#�B7#�̔"v��ƒ)?˳ea�8����]��
��rE���ƪϤ�Yk"1/Y#_Wӆ�q�©����0�w��ĲW��,)B�|aڧ������'Sea�8���`<4}��(����5�2���[@%����nEA�i�+���/?�s�m/C�H*�m��/2�ޅ���?�y��h��ؒ3����]ͧF���y: ��˘磋��w.V&��B֥�(����5�~���}҈b�-6F�s�%�}< V��,��B	hI�ˋ������Kp&�@���k���E����F�'n�^0op40�zɈ���y�,@���k��"�,�>E����\�v�)��+�}��]�.�b�;װ?�p��U��֜��3JHn��z����r>�L(\Ӧ�$�̎�)NC�lԇ�-{�v�ј�"��Z鎬���������o�	�7��r�=N�By3��<�]�!����M[��Ǣ&��s���q�����5	���]���>����CΌh��eZ�����E��@IE�U��>��l%i�-i��H�p�E����F7G#+��\w��0][�л���7"�,�>E����-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0/v�K7%'c��Et�p�VU��Jm�QA�Q* q�\E��0</���/�u��(�
t��Y�{'%s:3���5C�ݪ���CyW�f�tR�wX��hs�����n��0�5	x��(�
t��Y�{'%s�h�v���&���$S�ݪ���CyW�f�t<|����faՊJ�e:[e��mea�8���u�����B������"�k��зNË�����8��z{��E�EYZ/�矘��-n��I�?g�f��m�������d�k{��6i�^��s�n������9�3Ah	)ޟN���H݆�