��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�A���0>�kz��/ �_M��<-�[a�%�����'(�S��jS_�,��8��T�.B߫C|��N�(ݝ_l0fS!��mYԥQ��DF�S;���h/��9mϓo��ޗ���Fe� ����74p���D���<:\8���.��Jv�����%4�őba�Lltr��(�ubZ�d�m~�߼�I�&E�F��%4NV�η�fX���K�
��#d�
���s|7Ȧ*+���Ս��'1�U�>��CC�0��Z��l�+;Um3�����KH�8��Ԍ$ʣ��VjH�T_ |X�Y��bDR�2.,)�I�P��5`f1L���z��q�l�u����� �%�y�h����(�RP�q����>-���b0KT�$�}�� G��=(�g�,��G�z-���8�AD����}c��J�$��"C��Pvr���y.��D����a)gY������r��m7�l�8�)r�����@��Q�{8O��yR<q/��9y�R��,[n4C�'��#8e㶆*��jq��Z��,���q�d���R�����筳���o^h�R�<w�U�r7�b���i�"˪R|~l�����+�z��f�+���?9hZݸ���O��<sM�D~��b�%7/
C�]\���i.Z����z�:K�x�8�
�y{,�8'�3��QW�~ʮ"#޷��Լt��?�?9�	#(�s/v����
~�#%��I�}�C]v�E�G�R�`aշ�j���盘ۧ��w�����-��iV���B!Tf��f^H,��GSp���' 5�u�hB٤��Jx|I�z�a�sʏԅ/��Xd�_�Z��������c���쉣�|٫����)�E��"ѯ�&�|x/ݟ�%BQ�b/�)����+{�]9�=
�Cm�2SxG݈���֧�v�-�����	 �Ċ�)]a���)�D�?�����<�Uӳp�2�?m�&_x�߾|E�?Zf�`�7������D��QutEv��h��|�ӫ��:P�F㫉���U5`�/gz�` �fF��k��Q����V�;��S��ۭ��� u��bx<Ha\�U-X��O�LX�3oi��V�(b��G'_j�N�G�����(��fG����<6��(�;�����H�5w�B'�=���lq��~_8����|��{�Qj��~-���Ňz}��K&s�zzt�w�U�D�ܦ��gh�J��o.
���I���/�a�L�Ka���Q��_����؎27J!�p�	֏�
�����%-�%b����.�Z�c��pS��t��)��)��*���m�[�!��g-��HF�T�J�NɄ��	�D�!�t>r�3��[��b.|����q�&��8�U_9�I4 � ���B^_͖�g�����P��Ĕ]��<9�����U���\���ۍ1�Wd%6 ����;�6p[[5�*S�����{�0K[q�ۺ��L~�z���cI-���e�f�:���Dh�I/{T� a���ux��Z�y����8 �=�Ώjǔ~��������}����q7\f=	A��U+��q�G�i��Ѝ_)=���'DP�gM.e0��6{� ���o�K�`Z���A����3�Q}Ơ��e���#�7�Z������/ �=���s��.����*��e2q�<�O�!�qX��.��Ɂ�~/|�˶L$?o���g\����78�~�t�[�m��~8u�_a��1���+��e��K²T�q����ƭ��A3��."ïD����\?�Tn"���е73��"�u"��j>S�W�`��@N���2�1����D��q��^
��f� �P��wp: W3�H�TَIAu�N�C+�?����{�����ʼ�"w�--�>%�����6�)q�G禩ܯ�D�f��9,h_��\s�M�H�Ċ@y->�Q ���NRm$!�!Y��B�;�K>��o��ފu���ۍT�ZM��6��c���d��+	lIZ
�$Bu�`Ʈ���!�uQ���w��f��i3�qk��|e�'�¢�fXGe�'斋��g���}k�
�A��w�I�r�>+�>��#��v�aJ�	���y����M3�+x��	zj��"sF��=X�R�
�;T�R�'z��ە��%����*!Ђ�V��]Z����[������I�t��w�n%$;)�
�C}?_
�3��q]����\�|�Y"�U�)g,y�Fǵ�$'�̰�]�5����Z�#�D�=GF�´�j��G K*(a>u�è�(
��d��o�P&R!�?���Mn���2Q��\�y����֐��W�\p�|I!��G<	v[�L���_r�Aa=*E�X3�0�<B��DxLgyi��57q��U��Z��s��k@*�u�DY~��|����uV�\�oW������^�j�bQ�fC�\U��(�p�����W��cA湑�FCyX|���U�'(f~T%	���w����bQ�{l�l%k�7A�"������kD���������?1��}����p=�Ah��N��\B:�f��5�kyY��3��MJ�U�waOД��:m�!_G���_ѢO�����G�aZ�O%���A�'_-�Gr��|sDQ'������ܞ�*�w��U8��I�VP��z��+Oi~L��y�3��y�����ԑ��`ܔ�b� ��_4)I��Z연+�zֱ�d>.:BԖ���*..�u�D;����w+��C���b�Cq6>�/d=�5�;�U��dQu	�`��7�����״1��[<�u���}��|���L��e�T�m���"(m)���s�k��9���������۴�x�-)�6	j���y�odo�\=�]w�;:���+]EgB���PbZ��1��RU���n�ծ?%6Vm��^�ߵ;ϲ?~6]9@e?3&�o0��y��,id��^�@�����Ե�B�����E�i÷<*�#��vd�RN	m
ۧ9�m�+ſ�2�0cb�U�?k��-�9?�F>�Y�8�����]�s� 	- 6�5C���k"~�}�>�S2-ٷŀ�.6q���ޓ��ad�an�dK��~z]���H������	j&Wu�q=T2��Rt�۴*��$2����kգc��5��s��)C>���`�~������������N�{�x�-��f�ۆ��=�i�,D��2�?�}1�~Y-�/8�=�o\>O�v�L��=�jlc�����U�I�_l�9r&Xh>�su�P9����s'o��AЩg��g��N��v	IÎ��D_v�������� �dy�̖��aN���S�P ]K��ãS@K�J�͂W#����1�Kj�su3��V��Ƒ)՗��O�3�I
��6h)�o�����ㆽ�k�a͕me��*&�j�\X�e����	< ��5���	��T��Z{��r���Y�����w��r���ҶFV=�U�8��*vҹ��R���6�I��e���;�LtWyD�ov��1 ��r�AuCax]|�כ�,USV40�i�R<PM}��H�n�ے%���G�~�v��Z�o
]0K8�"5}o�"�݀s3��P#�N�AJ�����}�G�>8>�U+nNaM��d?�R�˩*��f���c��Wf������}X�5����w�Pf�o�Ц�IP�&�g���$�i����������5p�>��9P���>�u7zQq쥹z��wxUI4�iu���%�]cΊ����I����R�mN��e�͢?�A��d�����gC�C��C��yq�Z��c	u��I�����i0N�\�8c��ތR1siA]�{�ź9<��J�񞐂����1��'f�c�~]���y	 榤yw��yqx~��d�cy�K�,���iu?!^�ӽN��q"@�!m����G�� �L����[��=����\9�	[�M���&�.A��r�,m�w��䢍�=iN��*M�@�x@j�J��K�hs&�����d委{������Gj�i��Q�l����#/p�5pX7ޯ��F�$�1�|>(�n<�r�{p�/_7���5�>Խ:{�����r���Z��a���2?l�Ԙ���*[c���R*��l҃c�rO"}z�ڜ����6�\� ���XYj:�)ǿ�$�r#�TRX�XZ�^$$�֬0E%%jI��b�׫G3X�r�$|���6F3~�Wߥ^�&�r���y��M��3�C���9��צK�
S۷<�0K��~]^�^dw��q@�����������|bG���kQ��G���ѓR�EH��Oew똔�a�$�-x��P]@�`�K�J�p�a]4��7�7eq��Ґ��'�:&��»ǖ ڍ���p��r��@�*tu�Cʋx���b��3���k]T��*������ff= �t�ؐ��N����,6??}���֚7�k�^e��lIi�����Ϭ�[����φ�b�D��<x&;��4�+!���(�`� ��B�}��
�z���1�����0a�&&���l#�;��Ÿ#�E�F/o'���N�n�.�q�1Z��Hߔ�Ij��Ѫ�cHS&���@t��(Pe|��J����'�õ�<a���W`4?��n�f��
L�سZ�@��vU��2j�
�����oņ���n?�E�maPY� ���>�ʟ����I6M|!�VSԵ��f�O��Î��}B��)�Y��3�K�@�xԅ��{�o�G�\����� �ȥK��D��A�!�n�\Ni8��-Y�b��?/�����(,׆�,{m��`G<Yz�w� 5�Ŋʝ��8��GĊy�<D|�ǣ�A�Cc��� I}F4�Њ_�8��=U��"7-dA�Pe_B;����-���'嚘d
�yW4_�X��TJT�,�Nb�/�O���Fˊ&��0p��^�[ ._Z����G�C ��d`�d�oo�ȹ���K߃	���	�I�DM��t����\7������K>4=Ǭ����jq�o�*L��]��
�_n1F�=���ޜ�q�V"ڣ_��N\��R��饥�
%?� BD�%/u�5^�]�� N8�4G��S��_hH���vn����X�O�΍��:JR�H���p5�6r���@B[�1�f�bZΌ��iG!#|��q�`��19�W��kB�΋�i~�CƂ��{@��f��)�egEqz[5���$�v��%��H�R���Y�QC�x""l�S����0�
���y�����{���׿|آ�K֖�4^A��_>����Ah�ѧ���m"CLG
,��ۋj;��TeBJ�)4Ǒ��<pl�~&*RO���#�j*.v)\
/�X���&"����"Lر����������#>?f��E��aW������!����p��󺁽�ҍ�c����؀�<A�_�Nn����d�c�����L�t<U�4U����q��V�k�d���M}���� g:>Y,�vJ�Zz���g������!�0�S;QS�ղ"�˅l/�_-����J����� u�߮�$hK��2�7�0�C��s���Hx��@"bA5�Z����29Iwb�tH�.�Z�74��&�ĽȏZ��pZH�@!�����PE���v��ZgU0)� 6�i6��}\k7ևH�Ϝ�]��Ȉ���1���2�Ic�'�o�ЗT!Јt{�3zȱ}~B杏��ti\/�vj�fJ����ۋJ���6X��&��3	"ʪ�LJ�mr�Vx�px`j���I��-ʪ�YM#qA�=��d�����o�������be_��������kg�4���`2�V���g/h�O6�f���0
�����,��g�M����F{.�E�qZ�"R�x[�%K�n��"�b���P�\�&su��y���=�k��A?gꋠ����;���
� x�<�^��t���@F�I �D�ٶa#b�23�*h+Pw#�	��:ޒ�����%=�*q�' A���7`����")���@Dd� �)`+��Cm��L��g쭠��T����sJ�XQs���[u���b�b��[���o�o����kc�8b�������pr}m��wuB���C٦\���^+:%(�d���ª�k��vޖ��m�U���eG��D�����K�d��^��C,�@[=��o�l@�w��k��^|���y�6;6@@P<A�=~�e��� ��8ƟsH3�/��p�	�x	z��A�V�$��+Y�B��h� )>��=�wJ�͠�C��t1����g��#�΂�E�f� wK\z�=-A#7�D�������]�'J�4�@X�PF��&��\��^{�{3���l�������j1sy�kb��sR����oR����E���0c`� O��y��J��;������q��jT�1����DjY���Vy�T\?�0Bbs�� ���6�փ Yjۖ�U����;(�hx��=,�2�����_O�k��ֵ{س�MO�0���y���f���a3�(؁8eV�k�`�n�,8mi�SC���{����[;�ÂaybC�`o���$��Ac�9'��:���[>���'Y�͒�ȣ�>'
��ou�q/F27�r%���b�w��|4y���3�;h����M3��ɛ�@$(������TUA���wf��Z�NA7h��%�4�?7P(����g�B�X�ω2Z�Iv�㌊g^&�\ߵIiA�@x��e2�r�%�3�����@r�� i�wODЩi�e1HT�� O�J�d1E<��E7�;[�����m����(o2�
�2���Ǎ�l�yB�?8��F"\���i'���c��kP�����Z0m M6l� ��[[5i�%h"��30���)���s _��3K$��r����Is���{����B+�mC����kC+�Ϣ�P�`�������&W�=�bu�e�n#��������g��rܻȺ�sv�⨨gi
\��/����2�j&JE�ʩr�O�M�>5�H�?�6��A���W�
�6�ɓ�۔�J����R�AU���&mS1���W[��Z���Ŝߌ�[�?�r(�W@�n0�vI�� �g>�!���^��_�Qۉ`1-�%����r�si��e=�OG^q�Ps�1O�ȡ�"_�>��0����"��$~���qp�	b상��.��h����;s�$����X��X�~2��g��ME����^OUBBra���o�	ޚx'������vb.qM+����C�'̇�Y�����O�$T�ֿ���
P;�����]���X~Ė���t����[��t,�8��W6k$($�O;�U,��v�$/�I��tdf}s� �3X�ogR���h�¿Z����w�������^��&���gcTGZ<(���m!7`�V�mXՌv�80{�vY�w5	�K���	G��l����\B�
���rUkL:M�A�N�lG�]jY+��n�����?+R�`R_����S�X�d��z���H����/���hn\�5o���,7Z���zI^��e���z��K;N��Pyl����oX�+���p�� ���#1�z)��\��QZ�ב�y�匃�\�-,����NF��6�>���&K������⻫4n��t~>�GY٦o�Lv�}�4��H����
FJ;haI��,�gJ[e��+X#>`t������c܀;j�[Z�X���L��C�Uy�������gE}���R��^�6�Ӕi�w���#���:�(R*��r�I���
5���7�����!��F?��cp��r���<[�L9�J B�f[ B�����a���Li,�PGI�c��s'�e龶/ln��[C����:�%o�l��N}��-�o��#i#󊙸��uU���
d���_2��d���I��Z�2�ț���>lh�Έ<5�k�s#HHr��P�0��x���0���g>25zRz���<<�iƜ�4����6ͽj�7���I�Z�Ӄ�_���`u���q�Qa�^��k�,
Q�~Cz+ɹ��	�s�R�;\�����i�qX%��OyCy�6s�i*���Ǽ�+,��">��g�Ȧm)F�}��vlvB������������P��uԬ�/��M���w��Bq����O cB�~��W�7zD���d���Hm��X�\�����iؘ�`}��м���i��F��z��w�B�FU��$�����A��T�iQ7�=+�~��N���_��
�O�C$��QzOq9X߇�G��kV`x�W6%��x2y�?�D�y��7A=&�ҿ)ٽlJl�ad���7Ԯ%�<$�⺗���06�j�Ϟz���orL`DX���R���Ku�KKk/R�.T��[���71����ZA�]d�UTsX��(mU\<�7/�j �%���y�^�#w�/�h�X�9i��],Q���F���e��\�͌D���;����X�CLՈ���-��+}�9I9�<� ���R	�1�D�tU��[d ���{�H^�0��(�f��`L�L�dV�+�����a�-a�9�|�E�y�u��	&c��ƌ^�m�82D����5SRBL���(�8�0"��;�%����M*��p7?�A��e�d�i���p��0��Y%o��j��~6ZܚgZ+�qe��n.�t�@�H�J1#�_�:��ΉǦ�t)����P�����i�qc����f�5�P�1��"18�7�ϞQx�ZNl�*�yVRQ�?sئ�R�`g��y3GF�)ۑh���(�fv)T�zf8��$oK{��׻�{xVM�u����Am}i"�:/�i�u���<�܉GV,�$k�%�j���²t�A���5�a�a#7���!�a����[r��[R_��-C4Ƶ�ŕi�/��'���$��J����ʬ���X��������\Wb��[�9�8�\������/�G�K޲�kM��K싞�|�IՄޫ# �,Si�����y|�efG1p�:Uaѐ�vI4d�ȣ��l���4��1����1��{�Z��Q�3@6 �XM�d��͏R;��Q�9g_����{�q5���(�԰�������?�t��eD2K޷D��S&���Φ}�c��O�y��
Gug��p1�eW��8��I4����q��;	:��#0�v�ὑ+F�	 ��Dͮ5c�a��&���#<vN��[��L?Ȝh��?���IF�]���b��C˝?�k�DP���%�U�<���RT�g�>��c����~7n�����qt��Pt\
�e�!��r���ڞQrW�	]n'6�,�[K��Bt���୿��jbqD�Ϭ��Ac�>h�K��ע�ѥ���YF+�
\����<�ǡ ǃ!=nH}Rm\c��42t����><)� ��6@w�ȒڰY4��ͮ��v��߄�o$k(YX��؄j!*�Æ��ϝ��D�	�=(�fbp����dF���3�˝���M��E�5Ӡ�I#�_�\	���`��.�P�^GS�r[�>��R7��H0!5"t�':Q��k�]���y�������<ؾm������ �9�m�T��ylg����V���ؗP�	}�ஐ�f����o��r1^2�l�;	uD�%��P}�`f�Ns��ȩ|U�"ߣ�k.o|XXFs�L?�e9kN�tU��;�l�Zm�_����S�1�Z�X��L ���~�(�.�u'?E��ry�tj6�6Dp^P����1�C;Fr�T�P�ٿ87~�4Q1UT�8v�J X%�F˕K��W,'R�e�����&���Fc����0��~p�����|E��
�,5X��f�4�S�Ol)���f��}�z��nv@*��3E�C��9B��֢	�5!@7O�:��D,c/�	��IcnB~����.P���)��E⢙�u�6�(����3����N����2���SC)�R�7���(0LV5k�c�K�Sg�,o��y�S���W-�Įy���C&Ū��s�O5�	��-�dc���v-��`��1�^�0D����uC��5vw�ϫ�0�|澫40�(5�'
c#���ؤ�ū/�"�2F7�*�;�{�u�dA.��4�'aPR�7�C�.fzm1Nv���h�����<<�X��=�:�>Si�C1y;8i�t�f����^%+
���itrc�w� G�d�c8*f�	�pͣ�]���[ylj�?�:5Cu�s��5��c-���v;��k�f��ž8y�q]9ceIk-����v𹟺̰[�~a�˹�t����b�.S�<�3]{�T$��G>��K��90���(R~�w��e�	&l�'�x_���#����������7�k_19����:�y)u��Е�-�!@���m��'^���R�X�*����p I�*�����'�U�If /�Gr2�nKcC<���Z��[ ���>wC����p=av��%w�X:�����HJ�_�lvZN>�	�����g���vNd���ΰ9P��-�"�όr�+����?�!��ki�����f"��#��7	�e�(o�Nث�/tn8q����d(D}�֠�Y�����UDrh|�s�vox-^Y���1[9P�;��l���hጄ�åWEx�L��4c�L���o�](�h�n�#����
��U�/����]SR�����A��[v1'v� =�+����:I��&`��f�Mb��Tr�ݓ:Tqp)�$ВUqΐ��^�i��7��(�E0���"q�e��3����wB@�h
��M.�Z�� �5���`?����	��+H	�o���2B�p��/)���VFV��c�,vc[��jt��5�R<H�Qk���ۗ��x��끺	�U{?�Y���;(���:�O�9I�F�*��z�gpjȺ	,��735U���Ň�:E���B?(��<;���5I\��B3�RVغ����[�-��?��.�9$ �.�,�X�iX6`�	�SKW��'����[���ZL�f�����n+��"�Ш�-r�D���&�4=�Ԅ�Ͽ�7� �(���`}�kX*LJ���=��-�6�[K