��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����T�l䮱����<�2�]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPh2�ⴓ������g�ך��_�L���$�1�2m��+�<4��ˌ�ň��h������R��.�z,yN<��;��� B]�pE���	x]̃Dj#^Da����M�Ov��12È�pT�7y��z����)�,�˛D��w���旴4�����:��@���b���$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA��R����.���Zߧl4���0�?�1~�x�cK���}��P҉����D�YY�j=qvȏ�{<��t�����!/�~8���K������T&1h�9޳k�U�����ԗ|�*�	i!9�筎Ah��!�`�(i3,>O'����4�X#�Mwn���=R�E��O����&�<�Hԯ���Z���Jsȸ�"rR!�`�(i3��6����;g�(}e�$F�����` �b��0|]<w:��t��D)�\�aE+ʻ����o;�]��;f��H�h:qP�
]Ǥ����;a����+��퍤Vb�!�`�(i3!�`�(i3G����g.��{ֱ@��s��� ���G������T%Oc�l4`�	oO��z�8�]�e�!�`�(i3!�`�(i3FB���Շd�a^$���R�G��%��6�r���v��ʑF<������=6W����,@)=?��E����������m���
w<Y�"�c=м*�����iɐU��:�,-�r��b���Fz�!�`�(i3!�`�(i3��e��*�	�]��c �$d�I�v<�j��pW�қ�-��F4^���j\�����v8�!�`�(i3!�`�(i3�iz���<C �@nk�ꆂ�5�8�N�����I�_�k�8n�di�!�����Fz�!�`�(i3!�`�(i3�7>�����D/͘B����u(*/D�v�l�Ū�TD��荤>�k�����ׁgs�����!$B��$�.ni��l|�LH�F�m���,��~��P���^�������y�D-�Ur^Ҵ!�`�(i3!�`�(i3�����h�(=)7q�'er��.�޷��4���O�>�k}�r���ۑQEYx�q�;��{C��c�S+d�J�Г��f�u�����!-��B<ԧ�[��+��sȸ�"rR!�`�(i3�B�'��a�{�ç�o�����0����(R\֎u��� Sgȼ�sʫ|H�ͩ�QϿ�ey��<0!�`�(i3!�`�(i3����N����������(��K.�j��RB{?a� ~>>ը܅%Gbغ���:�9I�uEd�=�WT�%�i���*��W~�O�N����X����3�ok!�`�(i3!�`�(i3������!���C�/�y���ܴ�WM�P[��j�$�*7I���y�L�=sȸ�"rR!�`�(i3�2 /��u��
���ƸtU�����3�(�^��o�D24N<I8����\.Wֵ*&E�^8��xt��:_/�~8����A�߲wLB�w���#✲�@�킍�"�?���Fz�!�`�(i3!�`�(i3L�E��1I�OfUA`���B��ҙ����WH%���ܜ?n昼�2#:�^��R�8& .бx���cT&���@B�p0+�yg�ksD~O��U�Z9�P�P�q�90�_�'��'�ڭ�Q=^:�R���sȸ�"rR!�`�(i3�>=���#�	5��4�]t$;�o�O�jO�b�d�v:�ˍc{���sG̓�.WY��E��sȸ�"rR!�`�(i3�B�'��a��L,�X��4���Ʋ���CHbp��bxe��[�����D��AB�/A=��0����!�`�(i3!�`�(i3W]u�]a6Έ�%������+ך�^\DW}��Q��1��#^�����K��)F�Z�u6�0�4��3!�`�(i3!�`�(i37�s�v�ϿW�ܣq�h�ҫ'y]����r��>G�3����7�W�d@�����:߀�ׇӭ��!�`�(i3!�`�(i3��&�A\�M˩ֆz��o������(�I�?g�f���\X�<����8��U�[��Egܹ�e)�Op$=���uH�!���Ȗ��h�}�_0+��Zk ��U{����q_H�Э�LP�/�H
M��ވ�c�F�=o����"���	x]̍��;����k�7ꦍzlQXL����g&���ϙc�IK#���{��O��qC*�A�=#+����D�`5�vA�VG��M,������~�*g������_et�rZ�?ђ��P^(����gi���$R���b�>�oa.4��ۙ��x?�s�2zs���T�j�ߣR��zF�Y ��C���!�`�(i3=]A��O�T�`�[�����p:}�L���)	�8V�2�ԧ�fQX��G-�3��rD���Rb��Y�W�7��A�. �*rcxm�N�ɴ��~襊s�� �����p��� [�E� '���I����=��A]�;�J]�r4EG��L����~T�]/L!e*���e��)j��ӌ@�۰V��L { �6��}��%%��c�'GcoTAk�?������F`πѾ��/@��0e��H촼"g&�w)���Hѐ��tAa�/g�P�,-e�]Q��s,�~TM�e�w�G3�E��])v;P���i)���zռ��+��~��'���m�!=�y����h�}
�ԟ�dIQ�0^��-�:L�����Sd,�ϱ���	���Ģ/*0�(bq�� &@RfB�y�I[���b�/'��n9� �1�@tb��?�~���?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�@���rQik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW?���ʢG�M._�I�`D�V�U�'f�ٵ��xMB�9}��DG> �f�������7�����H�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR@�/-��E]o��in�m��+�<4��ˌ�ň��h������R��.�z,y�+(��<UC;6aJVlO/������V��r:O!�`�(i3=]A��O�T�`�[����
�XC߁���V�^�XI��o�E?
�gγʝ�Y՛T�QD�!�`�(i3>���'hZ*rw�w��Q� ~��
�gγʝ�w���f\PV��-�q����D	��U}c\(�T�m����1�p4/j��ㅑl��o�"�,�>E������m� �?�y�B���Q��v�[�D�v�l�Ū�TD����n̈́�����9���GAџVl��c��#
�NY���eb��D@f7�ܥ��2�NTګ'6�"ahD�G�bl��c��#
x�9#��#!�`�(i37�ܥ��2�NTګ'6�"��ؽ7$�	�s}��[�wH�HͶVq�|`kK��I����+�J������܇��cӄ�=�?�>��E&�|=�Í����>���'hZ*rw�w��Q� ~����.���!!?��~İ��K.�g�>���'hZ*rw�w��Q� ~����}2M�; �������@���k��l0��F��j�Ycs�$��Jl�y0[����	��N�Ae�#�k/�z�xEQ7Ê7�E�4'���Xw�������펎��{5��{l�f|�ό���.ӝ�\ Nhu '����'
���;���)"��%�����<��z��}�\w��0]vwdI���<�_�r�)�s�ި���`D��JU�Q܉zS�)37J*u>����CΎ�?����2�@No��u�Z鎬�������Ӊ*�@qO���o��C!T*�q���U��ݯ�AJ��=�O�<��z��}�\w��0]E]�tM1-�;��f 0�s&4�Ͽ8nЎz��j�Gn���ݤ>o�QݳwO�v��ՋM��y���[�ް�i".L
�^Z��|�ñ:Cx�o��C!T*Y�{'%s=ͱu���D�v�l�Ū�TD��������B���xBP��_c7�v�ԯ�'i�! ]���f�fx��V$�w�I�?g�f���\X�<����8��U�[��Egܹ�e)�Op$�jRE����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Pc,�w�&���#tvQ2�����\�w�Y��k��ı����;I7L���!��l8�������TI���*G���E[+���x��|T��j�"��!�����	Wm}�ȡ��b�2�k�%�w��6Y������SaB:�0Y�F�����#�
���N>�4�
��Ye�ήT�C�l/�8�h%g����R%iq	�g��w�?�b�>�4];ˍH��;[��癩I��'�J���3~�Mʆ�In��t!�`�(i3��xAE�g��Z��\_����*h7��k'�w��V�Ӕ�m�=]A��O�T�Pq������nk e��0�U�˰�X�R��%�������5���$�Qu��
Uc�v7��Q]� _�rs�i�����\��Ιa@�ߤu���.j��l�-��;��y�i����$�Qu�cT�Dg@�d�����rs�i�����\� H�ӹ��v�|[��N}�m��{A8�#�;:��MU��ԏ^���]/�"�~�26��\@�\��7s�9���o��S8�)qcA���_~��b�յ[+8�mxgQ�3\�Z��\_ՎKgkυ�H�RtV�^�D�����������w1���~H�%�swwI�e��+u8O�Ĭ	r6q�?����u��r��@�І�y��ˇ�h�͒	+E�5f	��
�Q�}������q�9�ͭe���PO�my$�N�N����j92�f��>8�0�������%!�`�(i3TaV*q��y� �ۮ��O�^d����Ě�����}Dq�f�d���yˑ ��Q�jR>Z鎬�������(���?�Rd�tŜ�}Dq�f��R'cf�����1y�N���kb�r!�`�(i3{�u1H3��p�.A��Vf�!�R,��1X�X�wو
	|�n�B�'��a��\>�R��ɕ�`UNP��ݓ�W���Ѹ�Z����4�0 L?ஹ�%�ԛ����C��ݚ�Н�(*�O�q(徥5B70�[}�N�`2���K���"��ӌ�r!�`�(i3E@�}n���&~e�e��E{��h����|�ј���|e"ʁ���Mյ^f�1Q�	Ղ�I8�y\��S��z�������I!�`�(i3U /숇�T�pc;�-�;S5b	��T�.,-���PF���6����3��^ؕ�U젩`#FW8�	��h����Ad���}Dq�f�G�&ց�*�n�sQPn���}���S.�3����Z��8�!�`�(i3pı��0��p�+^�ӄZ��3��w��\�W����-��"�ݓ�W����[DLk�g�4�0 L?ஹ�%����ͫ�CC�ݚ�Н�(*�O�q�Ե���[}�N�`2���K���)�gg>�!�`�(i3��� �C�&~e�e��E{��h
 ly�����|e"ʁ���MյU�K��<}�	Ղ�I8�y\��S��z�4��F9��!�`�(i3U /숇̹�������-�;S5b	��T�.��'�^�����6���u�N�,n��U젩`#FW8�	����z�&��}Dq�f�G�&ց�*�3ݣ/{�Qn���}���S.�3��ǰ7e �!�`�(i3pı��0����F�q�%�Z��3��w��\�W�Fd�.��ɶ�ݓ�W����߱v�`g4M�-S䨺ஹ�%�ԝ���,�ݚ�Н�(*�O�qe��0�U�[}�N�`2���K�����
���_���%>�rG�4���n����%>�rG�E`����y��j��k��0u�\k|d��1-���F��O�%sEW�o���開#c���܎�:��ɂHe�-�cݪ�i�<z!�`�(i37�ܥ��2��3Ù��i岦�%I^sb�d"L�i3�|)sՀ��UJZ_����>bL�'��Z鎬����5e �#H��6C Uؠ1����?��c_����+��O�IC­�4���O�>�k}�r���"X��[�~��yZ鎬�������(���Jbk-����'�\�n`��!��B�T�\ ��i3�|)sՀ�T:���V��'�Kխ�Bh����YW��b'�3Ai�+�t>�'���cEp	���>P�2-i_q?�y��t����k8O�M:R	�~��)#%�+� ��%�D�v�l�Ū�TD����>�֔،��t�h��W+��W�:�HCaIMl��ù:�h�=�	lK�M+P��˝Sz��E�4.@�7��y%%C�+߮��5˚2�<��B��ұ��E����.�g3Zv���� ��'G�+p�J��k�Nd�j��A��Di�HF9$��J��۝W~��0��w>��Y��$1&Od=��¾ȼ��Q�Y�+{���)��$x��M;���"�ٓC�KI[29T�y��S|�����,�A��N��Dk�_��g��V��*J k�oR2�����KN��W����E1�����
A�(H�]�z�	]��O5W!H�q�j�iT�s$Ħ��֠>�	�b���L��+�H��T -~,���Ho���da3@��[/��J=>���quA0�e]'\gWg��	�Z�kfcv�q21�ю��p�!-փ�`�5Ԍ������E����Fxy0�u��¤M�[�g��DW��ԅ1Qr�;�Ӊ;���eC2���9?C�ŧ2N��n�ܖ �&��ǳ<��C�
������:i.ߋg����$�Qu𙁚�^:�|�9��n�E5�����5	��)��8'���˟y�2N��n��ޜfbyQ���4��6�"y[�k	�I]�������a���~~]��Y�uߗN���g}�������\�vŜ�}Dq�f� ��b�FP&��㟷7��!�`�(i37�ܥ��2�'k��� �&�C�|检+�9�jɲ�1��� ����P�7� 1�ж� �4���܂��}Dq�f� ��b�FP&]���6d�!�`�(i3�I��?��\/ �m^'��D24N<I8����\.W��"X��[��Q[R�7�2N��n���ZS;��u�bv�N��y��bh��i�ԕ�j��2Vv8ۛ���a���	#�
�w��5����Ŷ�5YC�#�ڊ<?@U'(���d"����5'��èV\���F�`y6\�4�@�� �-j�1tSjv��]���`T�U2y�T�2'!�d�w251tSjv���6������S>��!�2r��	�sغ�#�/r�P!
�xI��P&�t�p�7�U�u�{�R�U�"7C�i����!F�G;��ɞ��/r�P!	"R��%2<�MF�~7�1d��]���M�敜�}Dq�f�5�����}Yms��/�u���4���O�>�k}�r�,0=]^	�&��|�B�����Yk��`
 ֢��؜J��vigܣ�k�g�G��X���5�p�mҷ}["��4���Iu���Jk| ǲ!�`�(i3�u��A�0���򴶽!`
 ֢��)�at��*��;@�1��/}�׏)#uE9�+��`
 ֢��s٪n�y��q��j��+��%>%��
�:qEp�;�P�t�5�B�'��a�Ƒ�^�2���B�>�G�Ro��>�������~���Eo^��6������S>��q�O�"pU���b��n��ELaԀ�8�}`V6�̎!�`�(i3�JO�'��`gw�T�с֜>�E�2w�f�%!�`�(i3/_�JIQ)vl.-���F1������$�����̪S�?-pm!9�>�:5A��p���F1������$����sR�I�uS+����:5A��po2p��8§��5<�w&`!�`�(i3�JO�'��+��K�L◁���*�8C��a������}Dq�f�1}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f�ϵ�֚��eL��O��pg��`�t3M)Q��Y���<�6�Q=�JO�'��`gw�T�с֜>�E�2w�f�%!�`�(i3��;kAbϗ���6�o����Ȋ�?ӳ4�;Ⓠ�X/�7�D(Q'׸��;�^�0�~�A���6������S>�y�-�RJ5Y�bv�N�ԑP�מ�����y��lDQ���jp���Yk��1}�ั):9��tf��!���i��L�p�z��+\��}Dq�f�1}�ั):9��tf��!��Ϗ�2�ed4���Ȝ�}Dq�f��1Ƈ��,���i������Ȋ�?ӳ4�;Ⓠ�X/�7�D(��S�����%��u����Ȋ�?ӳ4�;Ⓠޕ;j�j�������"�
�T�r�5��� л��
9̃Ւ/F��0��Jf���Ն� ��%�D�v�l�Ū�TD���7��y%%9���.:��Q?M8�f2;�jmT�#!r}<ﷹ�Q^�MY:T1�Ɓj9��jg����ΒՎ h.\���Z�
ʞ�^���@n�l�����[�ʞ�^�����t X��ݚ�Н�.$����0�*��D�x�=l�U�-kO��u�:�HCaIMl�i;��B��}Dq�f�`
 ֢��؜J��v�֋ڀ��'uE9�+��՝� s�#�BB�k���1��� �U��֜��3Vr�O���J�\���=-�aT����-�]�l�� r"�4EK�J;���[�uV?��?s�̵�7�!~u��r��!�`�(i3+ξ��?Ǳֺ�Z�6D��
(4��E2�DZ��w��뱐�!�`�(i3���F1������$�ӿ�F{ј�^�ݚ�Н��̢k����J�\���=��}��Y{Y����H�����1tSjv�!�`�(i3;Ε^����#��ߨ{���Γ8��������t����>PQ%cp��g�H���~��!�`�(i3E��\���Co7�wk���g�W����C�M��!�`�(i3����١�$�ݛ5�CNTף�[t�����������G�R�u��r��!�`�(i3AԢ�a\蟧��T�j�c�N��Ưb75���J>n]v1�_ُE2�DZ��[Z��.�~!�`�(i3a3@��[/�L��O��p�h].K��e)�W�=�k��:5A��pfĉ>99��A0ok����6������S>�y�-�RJ5Y�bv�N�ԑP�מ��
�:qEpCt�w#��@�ݚ�Н��j����D_���w�]Jq��BѲ�+���L>fĉ>99��A0ok�׹�G}:	�yW0�I��� 6q���V��	��y ��f"�`��H�A�ٗ��J�M�,!h�}�� �w˕�`UNP�!�Y��B
��v{�*�g!�`�(i3$H#Ö涅3�<_�ټ�G��z6!��Tޅiy:Vy�a���$�Qu�)�˥D@���f70���rA���oq��WX ��b�FP&/U��v&v��5�Ƣ6����7���~ֱ�q���Q��^��&sq�?��I�E����F�5F:	��ֱ�q���z�␥&sq�?��I�E����F�5F:	��ֱ�q�����Â�hfvL n9-�N�j�N�zg$�5F:	��ֱ�q��A:aJ�
Cj�R[zy"_�"tȇ_����ֱ�q�����m@Ǒ�5�o��7��E����F����o<rS�b�8Z���oگ��r���%��Q^�MY:��H<㕕ѿK��#�$����v���$�Qu�N�#f���C9*�¢ړN5Χ��F�,ؚ��XJbk-����'�\�n��6��	���`y���ֱ�q��e&-��Wn-�>[�@2Y��j�N�zg$�Z�>)��oz��KUq�2N��n���Ъ��4ސbv�N��y��bh��i�ԕ�j�a��ź����n4s1��7�癆cg��dc�@c�����h��-����m�0&�ܱ_��Nc�{ݞ�y��_��NcܦT�TN���s�Yls�<Ԍj��_�mS8<�n�ݚ�Н����B)e��0�|섃Va�ir�r���쳻�*9���-����!�`�(i3�R'cf��i�X!�!D��(J�f�x��2�+�T�\ ��[��(��!�`�(i3�]i �VB�۩�!���'�Ig�G{ݮƻ�@|�|����!�`�(i3��,!:�;��I,�D�y:#9�]�B�'j�j�Jy��Ww����x����VYc��M��̩�	g�x&�� q��j�J^!�`�(i3!r}<ﷹC����Խ�TЃ�Iʖ�袧H�RtV�^!�`�(i3�JO�'���)��B��YF�"���s}9_��Nc܆�v�9��!�`�(i31}�ั):9��tf��!r���ӓ7ed4���Ȝ�}Dq�f����%>�rGO�D mWN!�`�(i3�����$�D24N<I8����\.Wݍ���Q�Y�}!:��EM���
+����r�1��F���_1C�������9�_���1tSjv�!�`�(i3�gߝ�a��S\�$�8NS�p���]v1�_ُE2�DZ��[Z��.�~!�`�(i3`
 ֢��؜J��v�֋ڀ��'uE9�+��!�`�(i3t{�lPz��˝Sz��E�4.@��:u]R��GX�Z�X�W�NY���eb��D@fQ�ce�c��)=�,J�� ��C���Q�ce�c�Ԛ�-����!�`�(i3��r�Zw��}�@���_Db̟����O����ߎ�x��y�:5A��p!�`�(i3E��\���@cl��jU3����-X\!�`�(i3�̢k����J�\���=��}��Y{Y����H�����1tSjv�!�`�(i3|0u��\���.ޟ���T�E���U�6�'�)�Բc1����?��S(�`�ՙ!�`�(i3���Ȋ�?ӳ4�;Ⓠ��B�i.	���=MNԅ,+��}Dq�f�՝� s�#�K4ZRP�����9d��2���1���4X%��C_=A�H�RtV�^!�`�(i3AԢ�a\蟧��T�j�c�N��Ưb75���J>n]v1�_ُE2�DZ��[Z��.�~!�`�(i3`
 ֢��؜J��v<�8��k��vL n9-�N
�T�r�5�!�`�(i3���F��O��ݚ�Н��H�����7>�����D/͘B��< �b�V0e�{�W!�`�(i3���Ȋ�?�8�#�N���nJb�G ���)/��:5A��p
�:qEp'{w#/ B!�`�(i3�Cq�G������eV!�`�(i3�G��^��t��#u=�o�l�f�(���1��)��ݚ�Н�!�`�(i3E��\������Kū{rN���{��c� �o�X�!�`�(i3��Ě�����}Dq�f����%>�rGO�D mWN!�`�(i3fF�5.]����C�i��^!�`�(i3��~�lRJJbk-����>]��e�������T���ۇ�ݚ�Н����Ȋ�?�8�#�N���nJb�G ���)/��:5A��pfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�Z��/�Y�mr9�;ψ><��%K����`���t�T��?E-h���U���e��$�:]���\��5°ɨ�X�4�M�y�W�\/�ֱ�q���Q��^��&sq�?��Ijݭ�F���%,�������;���EWrqi}�Еi��os�z���+x�r�s�*�I�qcCl���<(���!����iE4���9�@�*8��ڊ��
��_w�7�rS��`���φ��<�6��R�~WI5�ZSV{:�xjzӝ���w3��׍�&�U��f�;�jmT�#�s��� P��#��s}������9�O��F�־^N��ܱ��*�������Ԁx숨�X�4�M��d"�S��k��'?"�ZB�!�_����^����ݚ�Н������]����o7��	ڊ��
��
��zq>�ݚ�Н��� �?CtY��zek�GHn�2�/Xw�e60���:]R"�Gn=n�k-�;��H`��!�fh����爮��J���ݚ�Н����F��O��;b�-�2��;�P�t�5�̢k���F�KD�Vr[/}>5��0�B� �b���H���������=6Ws��$�Z��-����;�jmT�#��"����G��Hb� h�ҩ��]���`T�P�|���5��t��/��IHy�Gj7�uzg�d�H�RtV�^;�jmT�#����n,��>]��e������Y��7����!�`�(i3<�6�Q=���y�� ӷ��ܜ?n昼�2#:爟yCje�l�B*�2���!��
`ϙb!�`�(i3��=�g�żפ	�?9Pjp������PN��7�v�ԯA��bu�x��ݚ�Н�!�`�(i3V	��V���$�w�d&i��f��`ȱ���}Dq�f�!�`�(i3�D=�-���@�.����ğ�.��RVP��m�`Őr��\���:=!�`�(i3.��J�ތ �D�q��E�b#�~9��c�	?�N����!�`�(i3���%>�rG�E`���!�`�(i3!�`�(i3~�`cC�4��.��cZ���+���L>!�`�(i3��'T���+��YJ~$��U:vĔx'�i�*ڃ݂S�����3�t�.K��ߎ�x��y����"ɻ!�`�(i3m|^�XlF��%�K�7�C��c�S+d�.�$z�Y�$]DT���l}s�G��P�p�{�MǓߥA\�M˩u���+�ʯ�`�D�ʆ�In��t��

2����C.�uE���h�/	��26h�W�5��|�����WāT���Aǂ<�'�/��YF�"����vz"Ȑ�7T�EXI����f_�������B!�`�(i3���W0�]��e|)0����n�=
�:qEp'{w#/ B!�`�(i31J\__m�q|�K_Na`wDlc!�`�(i3.��J�ތ �D�q��E�b#�~9��c�	?�N����!�`�(i3mv�%�3�]-�e��v��ʡ��
���,��;�b�0a*A&-�Ri!�`�(i3.��J�ތ �D�q��E�b#�~9��c�	?�N����!�`�(i3HN��R��Gu�"�0�!�`�(i35�����}Yms��/�u���4���O�>�k}�r�,0=]^	�&��|�B�����Yk��!�`�(i3T�8o��7�Wp��9B���@�ĵm�ݚ�Н�!�`�(i3���L2r{�"����N��Ưb7�Q�^8�bL�1p/-��N�]|-<P4T`�@���%�K�7�C��c�S+d�.�$z�Y�$]DT���l}s�G��P�p�{�MǓߥA\�M˩u���+�ʯ�`�D�ʆ�In��t��

2����C.�uE���h�/	��26h�W�5��|�����WāT���Aǂ<�'�/��YF�"����vz"Ȑ�7T�EXI����f_�������B!�`�(i3���W0�]��e|)0����n�=
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6��R�~WI5�d�֑���m/4@�s Oag��.M=��<�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h-�b�+�