��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���D7@aI|W�ϛ9�� ������[���a�8%`��4�s�6�XAoeuA�D3�O�þ�V��vMcr�|�zc`�G?q4%�}||�'�U��P&;m��Κ�P/�u����)O��Ξ4�"�\�� ���K�O�{�������>�U�۵}c\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\�]���џ�_�v%�]��4�:j�l�,9��I{��8�H4%�}|>���ؤ����2Ee�Y�R2
�I.��k��[/�!�`�(i3ئ�!G�?|lw��JF#�+�o���B!�`�(i3!�`�(i30�mv�a[�y!�3�'��sȸ�"rRQ@w�ӏ{2�����Vc2�����Vc?�٩o
Ή[Ed�+��J�+�2�����Vc!��.���jsȸ�"rRJ�a$�Y "+��<k�K��;`|/2�����Vc2�����VcN�RPLo�i��ԇl2�����Vc�aW���n����y��4��ʮ�:I��� %M��z'7!�	?�">�
Jf��t�c�.[K��m��ĭ]�	��B�j��h��UH&��?�ї��#)kP���{<��ha��׫��Dx�A�c���>��k3�ݑ�����Ic�"K$y"�hA	� ^��y�C���"���87ۺ�Y;����4��Y�jή-��8�#���@�v�>H@����A+B�e�u�阻u}�����!Q�a��*��&�Bz�$���ş@�t�k��V�W�a�{Z��h� c��(�U���% 9�6�'Mcö]mҢ�Y=�FD��}��b.3O�C�L���u��Z���a�\�nyU�-�Y@��#)kP����:p#e�C �@nk���0�r ��s���̴�uS4My$y}�'^'��|I%�&זds£����&����q�HS|6h.:;��<�..�4��N<��;���u��w)�S-!������~篟|�T��/%i���6�ЛL�џ�_�v%䆎�[�2N�8�#��q�)R������}Z�
d~g+#���e��k�8���҆�|n��I�� �U!Z���������ѕ�������ֈ:Y�x���' ����l��m�!=�y����h�}�Zn�h�+��>iG�ɹ�6wx���Sd,�ϱ�ϖe��!h~S܄=S��r��~��e������k�8���҆�|n��5�ɻ��Ͽ��b~�wf��Df����C���;���΅iG��w�վ~N���m�!=�y����h�}�~߈#���0�.�	�Z�@�@ OK.B����Ҩ�j�E���H�ٳ,�M(F�N��d�>�l;��r�O��C��0��?,*���S��I����)h�D��'����!�zg�Z�$�R�7��P4<�`�H�0�Is���H&�dcY��RL�a)�ƞ��U<��I��8�J59��Y<S#-*�)!�zg�Z�$H�2��p���:n##���Ψ�	�ǳ�V)WϷO��(a[�d����]	i}���~LɈW��^&�K9���v���y��֥2���~"VL�r��=1.	+��(F����"�����dhV��%C_L����c�.[K��mN,����0j Oag�?�4�ʗ
� �AH�T�t��3��e��ME
��偀6�=$��-�P\~KP��:�h|�m���rR|ӌ
r�����]B@�v��8b�m�!=�y����h�}Y��݅ 0�A�X"zB�j�ǒ��Sd,�ϱ�L���Qep��p�R��$���wT��xݣL��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ�^��+o���v'gn�]o��in�m��+�<4��ˌ�ň��h���T�%�/ң��Z���9&xc闑^����S��������Ǜ�>�xj7�ܥ��2��O�����ϊ���f��8���� +��u*K6HT�����Np�S��<#l=���E����F�'n�^0o��~+�ݗ���3^�����n����\�v�e�g����\Y�4Eb��Y{�o��eŭR±���]SBÀcۄT�٥��T����kF����K�ca�?��J��Z\�'n�^0oM�D�;��-e>����C8�����M�g����!�`�(i3��|g�Y�'���Xw��������lԇ�-{�Y%T��BPe.��xu	�>��l%i�-ʲ��U�4�E����F��j���0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6����^���m���>!�`�(i3c��Et��q���U��>�w�Y�#� ����������5	���]���>����C��"��K��~f�[c��Et��q���U���
��I��N�Cٺ�������5	���]���>����C�/$�ߺ��]�P���Qi��(�
t�ژq���U�[��N�������l�
H�w���]���>����C�pॻ}��!�`�(i3c��Et�Y�{'%s��.|Z���ǚr��y�_��wBW��8���/�y����\mע������Y%T��BPe.��xu	�>��l%i�-�Wv�4�1�>��Z{����|g�Y�'���Xw�j�7��a(􆿳����^��/Z�o��>��Z{�Ǖ�(�
t��Y�{'%s�ui�铨g��U-�e�,���6+����3rn��yn_Fu��TD��ό���.�>�Q�c6�`S��|���Yl���#�]�!����M[��Ǣļ$����"�,�>E���TD��ό���.�>�Q�c6곍�ٜ�]Yl���#�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳����^��2�0���Q�#<4^���(�
t��Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9���6�e�:r�"J��M+7EEN�p!!v*!����a0��\�ټ�]�����q���:�0a�0��+3ǆ/������}	���w��Ot+�z��7G#+��\w��0]�m��
��1���&���]2�y�Z鎬���������o�	�*ZV)�J����67G#+�Ǘ0z�cUL|�]���?.�9$[{^7��y%%\�HP@�a�~�7���� ��JL�N{a�9Ow�Y��k��ı����V���}���s+��� F���������R(��z�j�)�q��1�:�Ω�s8�R�	�}�����ֶ�#3�Ba�b�Z�l8�������dט�w��^���֮�LV����,JHn��z��p�Sg�3��ʹ�q�T�c�$�����2T�9�{uﱶ���_��a�\JS���Ux'��3�y_�IWYQ��)д���K�o�b��7f�R}�
�?�|� ���ܲ��+�J�����yg#��b!��u፠�w�`L�v�N�i����:��|}�
�?�pॻ}���'�gCm;�]�!��	Ǹ�y85��ٍ��%ڞN�gl��ܬa(􆿳���2����.�t������ֹ ��ˎ��U�g�q���U��@����gG9�'��A+OV��#��6�d�٣��v_���Zo��`c�N��nrm؊(�h}Nw���}p$_~R_kV\�헌�]�!����w�Հ�b02�O�uU�,r�-7s�9���o>��l%i�-5�e`��9�yݏ��&��Q]� _ό���.�}�
�?��J�'Ƕ.�6�G%&�˳͠m�xW��-#��k��b�`3E��Ҷ����PG��<h�6��R�A0^L:�b��tہpJ�f'���Xw�j�7���S�ڬ��M���q�tt�g��U-�e,%�0g���{.[��(�M���ٛ�~��`M��
Z鎬������_�,���R�A0^L��7rp��+�n`5�fK��0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6���2����.*X�Ɋ�m�
���n�)��X=�]�!��5����MW��)�`E5�Zg�x�ಠ�+�J��Y�{'%s�:�f~=g(���B���o��+eQ�s����|#9���b!��uፓ?L1��	���z�Ji��d�٣���N N�S��t�����}!�#�b����T[�Z鎬�������(�����-����28��m)a(􆿳���2����.�t�������V|C�ɍ�rH�ZZ鎬�����
!-�nlc��i��:�b��tIp�?�G'���Xw�j�7���S�ڬ��M���q�tt�g��U-�e,%�0g���z���Q���-j����O^3�T����0z�cULd�g>57<��ʹ�q�T�c�$�D�P�E6���2����.�t������:ux�����E����FZ鎬�����}�f������;�Ӏ��nrm؊(��@����gG�Jh��q-�y�� ��ϩ�]�!����w�Հ�*��9W���5)��Z^�n`5�fK���ġC���}�
�?� :b/�Ti��� L�>��ġC���p���G��9k�����a�|��_��^%Rx66ј`�B7d��n`5�fK�\w��0]b!��uፇN�*��	@"�,�>E���]�!����w�Հ�*��9W���O=�W�����+�J��Y�{'%s�ui�铨g��U-�e,%�0g����I��JnS��;	ȕ?���+�J���q���U��@����gG�j2��q�)��u�p+7s�9���o>��l%i�-��s=q�SbK����8-�����\Z鎬������_�,�9�+�\B~�S;��&�ˮ#��Gό���.�}�
�?�g�T�X�!�`�(i3JHn��z��ч��,1��;T��ኻ`Y�v��#s����4Z�1�#��d_%Ah�%4
>*"v%)��2��������� +h�xM��z�qg2�K?\�2�ϟP�зq8�Ј'���Xw���,D��2������ ��$���n`5�fK�\w��0]b!��u�V@���gx2"�,�>E���]�!���鉖�2ݓqE��6I&���#��1 bL�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc?��΃����7��Q*p_�ɬz!�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0M�|a)� ����35}jQ����4|��:
1�����I����~u[��l�,MXx�I����3rn��7�O�>4Bp'y����p�Ԩ����W� ��iE��G�����ٝY��e�s��6�(����m�(-	'e�F�o���^L�F�&�In���Hӯ�ɥ���؅��Θi��R#�K�|S�QQ5�:�b��t־u�t�6��7�L���:)_b���Ư�ճ�%�c��|[ht��p�Ê|��3�[�-aw�n��`�B7d��9�+��N�h�Gd��ނ�U�ɶ)g�YӅ:�ht��p���:�6 g��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�s�eШ,���	B8Q]D�	tf�2��I,nV�8,�y8n��z��t�b��M
rݓ�r�������7Î����RN�d?������lw��JF#�dnE��k~x�oe� 2Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha=�T;��W�.��A$�P������5d�	�+�&I(&�L��'ž1�|�'����u��r��'V`��b�TGaG��7Ů̢k���F�KD�Vr[/}>5��0�B� �b��7�wtMMV���W�I�M/*�3��E�i�m}6O�D mWN��ܐ�}�^�#Ҧ�����+C�!-lv0�9l{�R�$�V�fD��j��ٝB�q�g&�RΣ�*� ��o%���}�}ˇ�2F	��ًR���W�W�8�Y�
c) �1���!�`�(i3!�`�(i3]�xLW=9d�Ŀ��.��+1�����6k�إ��'�l\�=�]y������&���贵!�`�(i3��+�t2�l;���05�2��˅�S�J\7L��[����b@��)5�v��cg7Ԝ7(u��ݓ�W����'�ZE��ݚ�Н�����-Jg8�iT��*>������ ���Aؠe
�M����'����u��r��;�jmT�#�m���>#o�]�ʄ�v�4�?zmy�`��vN�[���}��W��L
�����xm�Olv0�9lo��l����� h�ҩ�9��n�7�Y���_j���(��2`���ݚ�Н��� л���:e �>���F*a��o���H�RtV�^<�6�Q=���ܚ��@��f�\%��WM�ڿ!�`�(i3��jVѭ@!�`�(i3�FW�DVx>74/��� �!O�Bl���%>�rGO�D mWN՝� s�#�=�U�u�íN=]8k��.ͥ�H�RtV�^���ܚ��@��f�\%`>��s����%>�rG�@�	����ʁ���Mյ�QP!Q� !�`�(i3��w�`L���ǚ����}Dq�f�}I�6���N�Cٺ��G��Hb� h�ҩ��H����D3w��'��b~*��s�l\�=�]y��d��-��!�"ǉ�t�����J�ϝ�5�v�z�7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j���(��2`���ݚ�Н��̢k��� :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3����-Jg8�iT��*��C�Y�\��Ra])n#Y�5�n����N6�������&G!�`�(i3VZ�ڋ���Y��<�{���
�:qEp�;�P�t�5
�:qEpj�E}4ظ�N�Cٺ��������� h�ҩ��H����lv0�9l�d9=���u��r��!�`�(i3��w�`L�P�~�9��}Dq�f��߆�p�h�Cd��9s��vr5�Dѯ���-����!�`�(i3�FW�DVx>74/����j����ʉ��%>�rGO�D mWN���%>�rG�@�	����ʁ���Mյ.&�K�F�!�`�(i3��w�`L�bP�[���˜�}Dq�f�}I�6���N�Cٺ��G��Hb� h�ҩ��H����D3w��'��b~*��s�l\�=�]y��d��-��!�"ǉ�t�����J�ϝ�5�v�z�7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j���(��2`���ݚ�Н��̢k��� :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3��V�v���� ���3�����&G!�`�(i3D�k���?���_j�����>�nE�ݚ�Н�9��n�7�Y���_j���(��2`���ݚ�Н��Ra])n#���r����!�`�(i3��w�`L���ǚ����}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3	���A��
�M����d9=���u��r��;�jmT�# :b/�Ti'ƃ�3�Y1tSjv�!�`�(i3����-Jg8�iT��*y_o�Yjfĉ>99��A0ok��fĉ>99��j���GpG�&ց�*�-�g�МQ�9��n�7�Y���_j�����>�nE�ݚ�Н��K�,ǆ�`�íN=]a��o���H�RtV�^pT/�GS�7s5kL�G��Hb� h�ҩ�9��n�7�Y���_j������
C�ݚ�Н��� л�1���~!�`�(i3 �4��s]Z�M/*�3�C#\�E:��ݚ�Н�$f��_Ub�F�S�1 ��̢k����0M�Ŷ斗���%�������&G!�`�(i36��J��c�� �����]M?��y�!�`�(i3���ܚ��@��f�\%`>��s�!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��!�`�(i3/�"����()�ƫ�w���>e�FW�DVx>74/���S�%�[KK�+��o���D����K�f�1tSjv�����l�� ��5%q���f�e�M?��y�!�`�(i3pT/�GS�7s5kL�G��Hb� h�ҩ�!�`�(i3����-Jg8�iT��*>������
�:qEp�gdq�_x�ֺq٫[�';��#j�ݚ�Н����y��lD!Yj<��[� F���E��a��@  ���@��w?����t^u�E�}ɬc��WN���&D$Aqm���W1!�`�(i3|����O�f�uǑc#˞�WT����Q1�'{�};�_�k�WSe��2LS#u�8�!�`�(i3���ܚ��@��f�\%o���LET!�`�(i3��Ě�����}Dq�f��߆�p�h� ��5%q���f�e�&�U��f�!�`�(i3��&E@wyT��$}�K5�F$��{;v����ݚ�Н�jCH�d*��=����h���7�)��~!�`�(i3���F��O��ݚ�Н����F��O��ݚ�Н��k��M�� ��F�����@�9��n�7�Y���_j�����9�x�\M�ݚ�Н�;�V&S�b�4���n��Fr��jL��[�)�jMOBn��akz�
1���;��x����2�K��n@�Xy|�W1F#�֞q&V��h���Y�-�:���0~�$ֲe���x���[��o}��a�lkEk=هF��[����n�/
�;�e!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�<Df��Eʨ�`N/��n��<f�:
�]�N������S�ݚ�Н�!�`�(i3}Y;�jn�����g.W�^�|��p�@OM.Ir�LL$����jVѭ@!�`�(i3��7I���Gf��x��9�k�n�=��M�{�|L���.0��AԢ�a\�2}$#h6��8{4����g��jVѭ@!�`�(i3��7I��٩h\K�5~�n�q�+�&Y��V����crצ��瑨R����q�ق��ӀS�B�.��iШ7^�	���r��  �fYCJd@!�-���a�.8�30�����a�į�vw�B��	���q��?d_�'7b7/�J�5����n�q�+��R�W�u�<�&�u7����pG`���IX0F�MV�ҁGG�.Mm-;�d=��¾ȼ\���F�`yx�>�+X�M?��yЃt����}�����9�lr�{��|e��0�U+�qbp@��Ra])n#���^a�nu4Bޗ��jw�	���|#HK��T�0T++�l��XulMd(ZDd�/��N�Cٺ���,k!��L :b/�Ti������s)l໶�,A/��M����,�,&�eǦ�@���Ԃ1*��ۦ��,:&Ȍ�g�F��6ð��T�ݚ�Н�pॻ}��$�2p[_��/X��-�����+Ut������F��O�}�	76�&�� Ӗ�t$�)�vxݳcF��kK�4+�ish�Ž��M�,!hޖ�A$�P������5d�	�+�&I(&�L��'ž1�|�'����u��r��;[�T���G�-�6�T�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����<Df��Eʨ�`N/��R��3���:
1���Ư����z���B� �b�Ъ���l���~#�W��'�Ё�')] q��j�J^s��Zf���R�o�"c�Pd�BR�~;�A*V�Q�� h�ҩ΄��������'|Fpॻ}��b	�fƏ!�`�(i31���~�����$λe�9�Č]2�lـ۞�[9o����HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}�-��cR�O�z�U����ؼQn!SQ�iʣLφ��<�6�@a� ��fFMqlg{y����i�q,?5q�I֬W.�M�4?�g�xjzӝ���I(͂��-����>�Q�c6�eK�	�$V�%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�<Df��Eʨ�`N/�<<��lpЙMǿI?���Y��E�܌��!���������l��[��o}q����]�+���J�2 z�P��	���QC�꠼*d�m�d��-��!�"ǉ�t������z��w3�_�]!�`�(i3@��	Ķ=�e���x���[��o}���h"`�{��b�b�*t��Ӎ���ݚ�Н��
�M��.��36T�.�[���}��4N�J�ף�[��hg׸��-�����d�tuѩT��Z|�F�̃��Hd�=ey+�8�Ȼ1��Rޡ�S)W�c�#6;8)
ߎ�>nQ\�9�	���
!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��D>�PW�� �[ٝA�x:��Tx��̢k����[�#��zuʖ3�z{φ��<�6��`䘸�|�x{^4��*m!�`�(i3���3rn<F�ڴd0��d����"��
��h�/�f��h��|��������aR�!�`�(i3���3rn<F�ڴdƍ2���l���Ě����E�i�m}6O�D mWN��ܐ�}�-��cR�O�ai��!hb�yaT��z��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���⛬]�OUbk�B�j�D� �*�Nw�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���
���q�89+�M�,!hޖ�A$�P������5d��n4s1�U��B��-� �ѕC?"�O=�W���7�癆cgQw�c4~Nr_�mS8<�nhDJ��3ZtgQ�9OZ����xO<�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b�Є�������O=�W��E�g�������(ӈ���m�r����6�>�@�	I\��Y� z�P��1tSjv���������O=�W����_r���9��D�y{~,�H�͛��߆�p�hج�a��Bަ.ȇ��_�mS8<�n�ݚ�Н��/Z�o���vP8i��l�_h1���d�xќ�}Dq�f����F%�᢯��0�Lm�<o��M?��y�!�`�(i37�UyR�j����^7����mgk�ԕe�p�x��;b�-�2�:䩒=]'HN��R���ء�I��߸��S�Ȍřy�m�����{Z$����}tM��楱�o��_�Rv�䩲$��8��I�:Fa�7��Ɨy�"c�t��t9������"sS<�0�zG�������&G�l�de����O|���/��kOT*qA����6\�4�@�� �-j�1tSjv� ���Aؠe
�M����d��-��!g��J�s��z�
1���;#o�]�ʄ�܃i�����'����u��r��J>zߋ��>ַ������?D�8����Ě�����}Dq�f�����,����0�|섃Va�ir[��l�,t���H[W?!\��쾇��i�AԢ�a\�2}$#h6��8{4����g��-��������C؆�1�u:�3u��b+}y[HN��R��bP�63Z�t�5ߧE4��Fr��j0C.�>��Vuq�/�Kκ~�Q��g�0��=�e
B%~��6�^�z�@��E��?J��W��x��[=�zɣ��S`&c�'N�jX���˫φ��<�6�@a� ��fFMqlg{y����i�q,?5q-�+���5wȏw�*��xjzӝ���I(͂��-������Ϟ4�>Ht�u�U%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<Dw\���I\��Y�W �+��}Dq�f�����,����0�|섃Va�irD3w��'��I�^$D���5i�a�vb�P����p��ݚ�Н�`&c�'N�j��O|������NM���$f��_Ub��7��G_���;�P�t�5�׹����忔8��;	ȕ?@�ߋ���|�G�me9x�a-J	�w���7Ἢ�i�q�&���`&c�'N�j�.T�Vَφ��<�6�@a� ��fFMqlg{y����i�q,?5q-�+���5U��F<�[F\���F�`yx�>�+X�M?��y�Dw\����ō܈��VW �+��!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^s�Uo���[;\v�a��ƍ2���l�}I�6���N�Cٺ��#o�]�ʄ�t�;��w��1F#�֞qj����#���:�I����Q؃�L�/�Ѿf���-�ྜྷ��H�RtV�^��v��7�t�K���m��"��ӌ�rHN��R��bP�63Z�t�5ߧE4��Fr��j������ō܈��VeX2����Ƥ��=(��9���Ih��t|��t[HNi�֌� I�'�`�_���&��"�*���"�k�&��3C��I�(�w}�tM��楱�o��_�Rv�䩲$��8��I�:Fa�7���⾰��bK���Ŷ�����\���F�`yx�>�+X�M?��yЈa�}�$�᢯��0����$�a/��kOT*qA����6\�4�@�� �-j�1tSjv�ըa��9�(�w}�W �+��}Dq�f�����,����0�|섃Va�irƦo�
�Ƴb~*��s�5i�a�vb����QY#��I2�8��[�@���=aS�H��ݚ�Н���U�R^p���P#n��뾦����%>�rGO�D mWN��Ě���aT��3G�IX0F�M�Uʮ�V(Y��a��R�%A���h; i�V�JD�IX0F�MV�ҁGG%4vkz����`���φ��<�6�c��:� �����"sS<�0�zG�������&G'9�и��{����@z\!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^����,����0�|섃Va�ir[��l�,t���H[W?M?��y�!�`�(i3��<�$Fo��<�����	G0��t�UW���.]��� 8w q��j�J^��!����E��=�f �T��ኻ`YJ�M����!�`�(i3,��B�K� |�>�
�:qEp'{w#/ B�t����}����**,n�4�G��rF���m¡HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}����f�M��-�5k\u�B!c�3Nφ��<�6�@a� ��fFMqlg{y����i�q,?5q�#���J�\���F�`yx�>�+X�M?��y��"�чE4�]�p� ��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#���N4�>y�pA��M?��y�!�`�(i3�ҹp3�Y(���27:�������&2��OY��~��<e�3�ݚ�Н�9O�m96��\��;�,�Ra])n#���r�����d�D���~�w�i��F���m¡HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}ĳm�����;}it�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��r�\��Y�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�9Ϲ{M�9�I�$� Xφ��<�6�@a� ���N��ȥ�n4s1��7�癆cgQw�c4~Nr_�mS8<�nQ'݀�=��Zg�x��/ ���we��0�U+�qbp@��S�!��EF9�0����ۏ�:��"��b+}y[4��f�i�Q2X��K���lr�{��|e��0�U+�qbp@��t����}���V|Cy�W�CbE��b+}y[�k��^�1��dc�@c�����h��-�����Jo���jk���%�8�Va�ir���+1�;�.��1���,:&Ȍ�g�F��6M?��y�!�`�(i3��QЪ��\��/���bx�F�{���!�`�(i3�?L1��	���z�Ji���M#�rYӗ��_�Írs��ʟ�r-�T-Ki�\�����Y,�֮����l�鵈R#�K�|TH��A>%�}שĭ{l�,��HN��R��bP�63Z�t�5ߧE4��\E�W��4b����A����q;�4�\����t�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��z��w���0��C�h�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcug7N�RL��{��� φ��<�6�@a� ��fFMqlg��èVxjzӝ���I(͂��-�����9lD��XH�|ը�K�QdN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�D'm�����Z<��A!�!*��*8�N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s��ݚ�Н����V[���*φ�\-�gM�?L}�7�n��<f��5p�T����՗fc<1tSjv�K��ft���-:��;��ч4H��&��;�T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH�|ը�K�Q5����{�q��Ɨs$f��_Ub��7��G_���;�P�t�5�׹�y���3w�9�ᾓ'�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!$W�j v�'���H}�@v���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h;�ƽ�/����zN�S���t�T��?E-h��`f���sd=��¾ȼ\���F�`yx�>�+X�M?��y�P#+_]ݱ�m�
���nGW�:!�E�/��kOT*qA����6\�4�@�� �-j�1tSjv�X19�-.|}�ڎC�?�x��w�����ԬQ����5��t�	���QC�꠼*d�m�d��-��!|�|�����@��pr��4N�J�ף�<Jq�Z9�`u0�F��a�Va�ir�À���<��aEG���B� �b�ПB�'��a���{y�mV8��0��1�"�"��K�w(T"c!s��̢k���
�I�8����q �H�%��ZtV1{,�m�ښ�-����P#+_]ݱ�m�
���nGW�:!�EҰ�WDChFb�Ht�!fĉ>99��A0ok�����F��O�\E�W��4b׏������{y�mV8�	՚�^��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������]މ�;�Gۍq��e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!@+�ϕ���q��B�`�J�ɉ�z=� ���ɡgJ��E&(p�
�Eu�J�?Ig�(��9��ᩃ	tN�\c�-2���S&ϊ�;ѩ�E��p��u��.t�=EpH��j��A�0: ��q����%	�3)���C*4��]���
@�i��g�?�d���&�V��o5]�:�b��t.�C��6�o8:4ښ�*jl���C>��ӚH�RtV�^����Y�z0=�_���{_8�Y��=�}�Vݨ��}Dq�f��R'cf��>��YfG��-}RY
xǍ�J�r��ps��u1,����Uh1�[��(��;�jmT�#PB��/���߰�$|�Pu��r��;�jmT�#��	�DůI�߷�c/��-����!�`�(i3Jº�FO"V'PS�����S�ڬ��M�kDu�H��Ⱥ�Q���'g`$�YD ��� ��?D�8�鉅�%>�rGO�D mWN՝� s�#���k$ �H����ڻ�+���i��ċ�!1tSjv�!�`�(i3
/���p\"�!˥���KS����<;�$��\|����=�'�^�����ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ��?�JY�)�,�Ջ ��C$�)�vxZ`�b�0P!6j�"Hsކl9�p��e޸XhZ]<�����	��TtU��
g1�MVjg[؎��&���.ԥZs33� �=X����\�5�O�%E#P'}�\$I�}!�#�bM�,!h�z���#A�}?ɝ͇@���8-|�D�7��aM*:�b��t�l��p�xB�my$�N��o�/���;�SENan&�� ���� �KS���*�oF���cԱn�+|�[Xs�g��������:=�)��S�2�]�Q$iP����p��ݚ�Н�X19�-.|}��FL��G��Hb� h�ҩι�+�t2�c�^[v�5�ܾ��mk�9$[{^+#y��MxOܳ����|e"fĉ>99��A0ok�Ra])n#���r�����Jo���j� ��7P��'����u��r��!�`�(i3����Y̀�3#O�2�B���s�����X�X���`��,n��뾦�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�fF�5.]���E�i�m}6߸��S�Ȍ��9�ڮW;��|Bΐߧ �l�}!�#�b�$2j�K_ryQ�j6�S�z�����F�t�ϛ�c�.[K��mZ�'����Z�G�a}C��B�No
/���p�U�.��k��~��/6�o8:4�I���c�90��G��6�(&�L��'ž1�|�'����u��r��;�ƽ�/��e޸XhZ����xO<�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H����D3w��'��b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z���܌��!���uxrBZ@2`u0�F��ay�z�v�À����@���l��[���}��M�?L}�7;Ȼs���ݚ�Н��T1�8K��}!�#�b:��c&<:�b��t�����W��k��^�1��[��o}��MX�w����D����K�f�1tSjv�K��ft��;�cM���/.�,/j��O�`�mp8V��%�TgR'��}Dq�f��5ߧE4��mJ�0�6�$f��_Ub���uQL+��φ��<�6�
/���p�U�.��eWo�A2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܺ����ܟgx�/.ؘ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������c����}�I��}ܚփ�c���A�N��'���#����x��_�ΙB5��~�6�o8:4ښ�*jl���d=��¾ȼ��C7}n���R�E�g�������(ӈ���m�r�����i7N�_�Ar��� ��w�K��ݑ�][H�#Sv�Dr3�'g`$�YO\����*A&-�Ri�)��S�2�]�Q$i��a��ݚ�Н�����SP��'�K �_�mS8<�n�ݚ�Н� b��tY�0�����V	���Ċ��NM����Ra])n#���r������C7}n���R����c�Q0��b+}y[���%>�rGO�D mWNHN��R��bP�63Z�tfF�5.]��aT��3G�IX0F�M���3�#<�W�'�B��"Iե�䛑��e���kn%���-j����O�ct���|��U��'"!�U��)���Y;e�iK!���d.���+�^n=\f�5>�� U�c�pl�Ф�T���r$ɓǃl[�Ƶ�1tSjv��m��
��>W�~���%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�m���>#o�]�ʄ�M��,����q���f�e�x��w����֯���,mk��L��q���3�tޙp���/�dI{�n�|�-3��e��2
-�XC�������,:&Ȍ�g�F��6�2d�I����ݚ�Н��W� ��iE��h�{:m�vW(�����C�Y�\�T+���f��,�,&��`�2,�!���������d9=���u��r��9lD��XH�H�߳Mk��{	�*Nx����O�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�]~j�wҍ���]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�`c�N여��;�Ӏ�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0�]y�Q�'��3#2Ex��D{��#!��׏��Z�׽i+�ȕW��L
��^օ?D^��MQ���0f�Ϡ�����b+}y[MQ���0�-��h���i!��6j�"Hs^�Z�cY�Z��~`a�K��j��A왏3#2Ex��D{��F���ˏ��Z��C#/<���q6 fd�i��sM}�!>m�Z9a\�-eO��v��èb|5�;l������Q"}Hi��v����o�A�,�
=���f�,�k]�c�jd�L�N��Ưb75���J>n�	G0��t�UW���.@�n������O%��}|�[]?=���N���9����v���V������yآ�D�����尠"������d�bv�h�C��p�@OM.Ir�m���>#o�]�ʄ�M��,����q���f�e�j�5˺����D���.���z�<,�\δ!�}�fb���l!c�ڀAԢ�a\�2}$#h6�ćm'_��Mw#�vzR5�<���X��O���r����!�`�(i3�>d�g�KR���8��h�	�O�zφ��<�6�@a� ��fFMqlgd=��¾ȼ;�jmT�#bs��2[�a��o���H�RtV�^MQ���0�-��h��ƍ2���l��k��^�1��dc�@c�����h��-����<�6�Q=�y'��BS�6n��e�<y�������H ^muN��A`	`#&�Z��1�O?rof�B�
�о�J<������j��H�߶:�3���.�BU�h����;��#�a�Ą�����kO�d��-��!$�)�vx�;�U4�I�';��#j�ݚ�Н���f�,�k]Cw�Hm��/��kOT�Ra])n#�ґ`�g�y z�P��	���QC�íN=]b~*��s��ݚ�Н����a�so!�}�fb���l!c�ڀAԢ�a\�2}$#h6�ćm'_��Mw#�vzR5�<��KɸǑ��)��#���?{����;�.����^����>=���#u��r���#�-�p�G�6�!~�n��뾦�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j�@�f�smy=$o��ɝ1��,Ƌ��6j�"Hs#�{'�?~o_���B䁒_[�FquA0�e]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7�p���"Fi���*	\���F�`yx�>�+X�M?��y��#�-�p�%��a�����b+}y[�k��^�1��dc�@c�����h��-������#�a�Ą/�dI{�b~*��s��0M�Ŷ�Eʨ�`N/��R��3���:
1���Ư����z����-�����#�-�p�%��a����"��ӌ�rHN��R��bP�63Z�t��m�5h1���g�F��6&�U��f�!�`�(i3b�6��R%��v�ډ��%>�rGO�D mWN��Ě���aT��3G�IX0F�MY�J+�WTI�;}it�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc4�`�(H��L����M�,!hޖ�A$�P������5d��n4s1�U��B��-_S���\��uW������r$ɓǃl[�Ƶ�1tSjv�t�R!ME�'�^��������@|����^a�nu4Bޗ��jw�	���|#HK���4Y{]$�AՁ_�mS8<�n�ݚ�Н���Q7lY��)P<�ܓ�Yfĉ>99��A0ok�����F��O�\E�W��4b����A�ձ^�Qb�Upq���!���_2��VU(��z�j�Aa�R�