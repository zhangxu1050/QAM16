��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�*���g S�ĲW��,)�]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPy�����h���!�}�1�:�Ω�*���g S�ĲW��,)�]P*m����)O��Ξ4�"�\�� ���K�O�{�������>�U�۵}c\֣�I��B���t��|U|�/֚W����͇M��Zw�U�;�\��"O��Ą��J��]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�Kwz��
����J��$mm4rz��x�@@m	G��{cB�38���E���2O��'HY-�������D���J7"-ǋ 4�i� ���������	x]�<���eQ���X��\���|�@c���Կ�:�%n��e�ι̕��R)U�~�O���`Y�5���=�zX4P?�o��ľ��UW��͌Tfu��w)�S �J���vy7��Mv�9�h�s����b�z�Y8�:r&@�	��Ϸ)�����V\~{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�T�`�7?�\��4�/�I����D;�~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/�R����+��T��M��j@�����nEA��Xc�>г�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcJe`xҖ3Ӫ�1?)�Cu��şo��q����R�_8�%���7���%%�xg��ۺ�D�U���&��,� A���W�F�ݸ��]ds�lOLH����DK�$s��?xA4��?�d���&�p�m~|�֟j��?q��N���%�5<{��T�O���6���\q��+��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc'.O��m2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h9��)�N6mj�N?����;t>
S;c+�«���A�3�+��Pŧ|��aN�A%iߘ�kKn*i��5>$c��8��-��+8{�7�D�`����)��o|�S���w���_���`�?�b�����[A?H��Z�!
���>X�J H��K�zk�����x<Ep�����Beba�O�P�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDLY�m��?H�(���B��������
��s�����E���%�a��s�����́+N�[�I�AJ�㗲F`�ю龀�k"Ty�,tT��A��蠿����d�Uf룘�_�]�|k�H�!R$�W��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�!�hM�-� ���]����;t>
S;c+�«���A�3�+��Pŧ|��aN�A%iߘ�kKêM�.Ze����`w�=�ֳ��ϟl9�ղa?�x���XT�G�*J
1H�
��M�� O��:}�w�?�b�>�:��^L]�'1�w�z���vL�vO��Ej
/p4��?i�������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開Ht7s��֨M��n������B��!�>��y�3əLܒ�� H�j�(A2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��M(?^v����"��y���D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���[���RdM�5���&��X��#����{�N>�4�
����`����������
%iq	�g��w�?�b�>��]�!��11<�InN:L:dK}g\�溂�;�}	�ф�QSg`�q UT���u�I7.���K���xc�1������
%iq	�g�须<+���UIK�tđ�I��U�;��r O��M&Fo�����X����t���skJ�t!$4vHv�߼
�d���f�����n��i���F�!�� <&�M#�4���7Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���6�x�%C��m�o�GŌxy�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�;����-���i�L��$�t��LF�E'���q߼
�dU3�(��M������
��8���i��,��a�8�
,FIݹo��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc?Gu<��\U�����z�j�P0�.Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hH�*)iM]��s,�ӡ	��u���������`9k�aa2��A�-(�ᦣf�߼
�d;�"�7� ��5}�Y7s�9���o��S8��@糺뾃7܌:�\w��0]߼
�d;�"�7� ��5}�Yq��T��h��<�q��7܌:���ġC���H�*)iM�;<XD������p!���?cC��O�-w��^l���Q�>4�b����"��y|�
�xr�ȳh�L>s�]�!��	Ǹ�y85�E���%�aS�)37J*u����k���開-�J4p'�>��\��:��AԢ�a\�w�?�b�>��]�!��11<�InN�Sc�j H����/�ʹ�z�$�W�@��!���~Pw-�h���&��t�F߼
�d��5B�!d_�4�yQ��o2C�g�kgw�"��I66�v��Gߕ�bȃ�J�����ݫ�����xoϼZ'��io��w�gӨ*Y���wYDK��R&��LN>�4�
���o��QNj�4�yQ��o2C�g�kgw�"��I66�v��Gߕ�bȃ�J�����ݫ���U�"͓�<Qs�$ʧ�x��S&ϊG�mU	���T���u�I�Gl�ĵX�Fʪ�t�����D����q7�F �Sup�xg�?�qi��g4;��K�γ�:�K+`T���u�I�CR��Ի��]��I���DƯu&7���F�!��t��\����b~�ff7w��fы��ξ\��q��C缜�(���Śę���	`�H���+��䓿槶q��T��h��<�q�`дȣM�lr?j����è��rTW|xڽM���t�� ���OgۈPM�����8�}$|~ïSup�xg�?�qi�N>�4�
��Ʊ���0
rcLd̓��>8��D��I�d�X�VM�����a�"�_�����Ӫ�W�F�R��
�=�1�:�Ω�*���g S�ĲW��,)K0�;����"�|�E+��T��M��j@�����nEA9&xc闑^���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��	���X��a=tY"0�a�"����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDLY�m��?H�(���B��������
��s�����E���%�a��s������XP��~�26��\�o�mW���5F:	����n4s1�ЂDa��(�_�R�G��=�gw�⽒��Շ9�/�|#HK��ehj�t�����U��+��-�����y��j��kQ�gE\�;��}Dq�f��5ߧE4��HN��R���מu��� �H�0��
�y�"�V��5M��z�o�:�Jr0���W㇪2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���(���c�0C�n�j{	�	Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y�R���1x�]�^�[��n��iܕ����������a�"�Z�>)��hC$?���;���EWrn6~��c[�3C���_�����8-|�Dp��xs�S��\��;�,�i7N�_eE
��'�Zgt�n����H�����T6�<��+H���3�u��r��Ƹv��*Qx{mw}G�e���%>�rGO�D mWN�u��A�0�Ή*��a��t���
��{�<Ti�2��-����Ƹv��*Qx��~+�ݗ��Ě������������0u�\k|aT��3G��w�K��L�V���Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �_d�Jq/W��]���mn�j{	�	Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��C�<w��>�8���Ę-ai.���@��8���i�E̳&k����_/�A"�U���w�c*����N��N�.`�Z�����èV$ Hl�]���'�PD��R'cf���_ľFW[��(���Zj���
Ӷ1���+H���3�u��r��Ƹv��*Qx�*��,6
�HN��R��bP�63Z�tfF�5.]����C�i��^ʥ�nr]�b�N���u��A�0�"Wm��|�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-�����!�HAv�r�G2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��yu��fD�پ�n��i���F�!�� <&�M#'���Xw��`UNP� ��b�FP&���P��'���Xw�8&���I���|I�����ï��9_��z#��#��\�Ж ���-3�s�T�cΘ�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��U(a��,��D��d�`^�ǈ˦lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL@
H$��jg��+˘\5;ԉR���Fȵ�ixUS���<+���U�"5� �S�֯.I�ұ%iq	�g�镘`UNP� ��b�FP&���P�����B7HSSV7�pB�R�wX��d=��¾ȼ;�jmT�#�R�\<۳��Z�^��� K�bXox�!�`�(i3�0\� ��+�R�\<۳�H��ׂ!0��ߪM3��J�g[j�"G���b���6DI*G�"rs��{|�����]�w9"x1Z���
�;b�-�2��;�P�t�5��=�g���>��i)�'a>-#�}�7��[��(��o|���P��3 �n�R�]c�����u^��󀋄�g�?�JY�)�Y`��jD4ЂDa��(W)5S�7KnZm`�x����Cҷ��e��߬}u1ʥ�nr]�W,�9�9<��U��g��+˘\5��B�1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�<	)}(���۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d���f���:�t1�$8h��<�q��Ӆ�)�o�A���l�N}�m��{B���T�D�a�x��nק��׬��vGC���Q[R�7��èV$ Hl�]�ǚv�j�3,yĦ58x_N9=rE'OR�@�6�֐<b��5^,���qS��z�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����R䞿�K�R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��ш~���}���i��ܕ����������a�"}�=Ll���]�B���[�^����[Oa�k�],��׼���δ�C[�����ͮ�px�����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vct��C��w�x썅J�f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX��"nq���z_�3���4�듴,`Y�{'%sa�6���� <&�M#'���Xw��`UNP� ��b�FP&���P��'���Xw�8&���I���|I��a�ѨbRi���Qu���%��,�,
((�H*�iH��[��(��Ƹv��*Qx�2級|(+bc�ɾ:$r�t�}iCt�w#��@��S��c��څH�8��)B�>T���u�I�F�M7�,ޫ�^���D����q7�F ��W�A#p�VU��JhC$?���;���EWr����Ly�Řq���U���n4s1�ЂDa��(�����U��V5+��:�Ąk��m%�l|���*A&-�Rip��xs�S��L��F�g:_���}��E�i�m}6�E`���ʥ�nr]�b�N����LE�Z�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Jl�D�&�/e���,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I��U��؀N�&jl�o2C�g�kgw�"��I��R� V�pFr����A"�U���w�c*����W"��ό���.�d=��¾ȼƸv��*Qxm�QA�Q* 5�����}Y�]��h@�YyZ��}�Q?M8�f2$ Hl�]���P��))O���w�_fHN��R��Gu�"�0�R�@�6�֐����o��4q�I�w�o���"��y|�
�xr�ȳh�L>s�]�!��	Ǹ�y85�E���%�aS�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3���/��kOT�i7N�_	�z�w.{��w�_��(�6k�4d�{j��b�ڐ]���!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���QV��W�
`���]{s-@Q<���2�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vch��\��f�U���e[�.��<PMאI�|��;�+ɣi�D����H�xd����)|C29)������JE'$Io��Zy��iȱ�K@���%����J�$�d��d�nĖP�j��D����'4ꛤ).�޽���F~h�����"��y��!���~�Z27B>q��T��h��<�q�P}��O��ꅽ52�����8-|�D��=�g���>��8��-�Ϡ���:=T�zU�k�I�߷�c/��-�����y��j��ky@�KF$��}Dq�f��5ߧE4��HN��R��Gu�"�0�R�@�6�֐���,���z��V1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>���;��4�h�R��4��N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���-��ԣ����/�ʹ�z�$�W�@U7��@��5��<�>��O�J�l���d�-}L��x�kk8/H�T_(Z6����g�q����h~S܄=lx�����bLVuA��h�#� ���Jp�1jN>�4�
���o��QNj�4�yQ��o2C�g�kgw�"��I66�v��G���V>�R<d=��¾ȼ5�����}Y��	}�@��`-z����:N�:�לQ?M8�f2���u��o�t]`!�ð��T�ݚ�Н�6�����l,��HN��R��bP�63Z�tfF�5.]���������G�}:�$B�>�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�s��rϽ��<T她o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڲ2ꧧ��*�U�"͓�<Qs�$ʧ�xX�,4�?n.1��ܐW�܎a�I���開���ۆ�#C�2���_�	P"G�wk��a�S.l"��<�W�C%���6V���~�26��\� :����jݭ�F����μ<�e<�l��Tc����omi7x�	��|N�`,9�H�Wq جI��A����� ���	�|���H����y(U���������u��r��uD�*'��'��{��I��`j���%>�rGO�D mWN�u��A�0���򴶽!��pM�J�8��`��4q�I�w�o2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �����.��cr剄u�R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��F��iW[�`����C}���D����q7�F �}x���cܐk�a�A"�U���w�c*��s
�%e�4�v�{o����
u��8&���IS�T"�IÉ��,�,
((�H*�iH��[��(��o|���P��3 �n�R�]�sN�D���l���}�	76�&�R�V�"�0ɶ37y������(�;-��LE�ZKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h?���ϙ��(��9�M��N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開I�	�*����D����F�r�m�3�37y�������x�W8�{�����!�`�(i3���y��lD�y?��as��6���n6�<|������`UNP� ��b�FP&�����c��b�Bϱ�{��<IĊ�g��U-�e�{g�w-��-��/$�i7N�_	�z�w.{��w�_��(�6k�4d�#��M&s��_�?<��!�w(�y?�?�JY�)�֬w�J%�H�V�®zz ���-3���<Prt���o�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��6n-��a=tY"0��N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開_9�R�5;(38�b�Dȼ�\�v�w�?�b�>޼�\�vŕ�`UNP� ��b�FP&�5�+�N��B�)Yd=��¾ȼ�Jo���jN#C������S���*�y��j��k��%&�gN���F^��	��x�(�6k�4de��S�Ò��X��{a����F��O���S��c��<ך{�X���/z*x�n0u���g}e.+�Re72�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�������{Q!X?[��둞���]D�@��z2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�j�P�tCu^(򎍖=b�b9���D��8�硤d�X�VM�����a�"�'n�^0ohC$?���;���EWr��uNS\IÙ=�H^����zj��èVxjzӝ��$��C��1tSjv�p��xs�S��O߅�Y�E�i�m}6O�D mWNR�@�6�֐����o���X�#�T����o����S6]Z����>ZB��}�I�?g�f{ì(Q[nS5H�j.F�6��^��