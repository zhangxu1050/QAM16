��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>c��mW���rJ(���/	���~J`2F�x���4W�0V�y��l]��X���8D�G$�ۻ��c��rk�E8o��W��z�����O�Q�F��?-_�䰹��Ny����o��:���l�,�:^�G���G��ta�`����k�8L�@�!Q�,��E�E��_��2���)ֈG 9X?#�ʡ�7��	�g
>|����.-=���D���I~j�y��EU�K6"�����=Tؖ��.r_�6��[�q�l�˿�B#��0#L��#T(���X ���Z�L�!Ց��f=�B�П�ī@c��zV	.Zp�d��p�3�[H�P|�p� �_9�q8��ژ�)�ƹ�L�(�p ?c��$���y"K4����~��NZGx�����(��=���8��Dѳ ����!�aPiW�!�[�$2g̏���Z�g�OS�o=1�j���ӡllc�:P��j�Ls�'���8��_cF�4�������O3^em�U�6cju�-v��#s��~ev�f%qNL&���>�,� gyQ�"����o ��b��}%�u��aPy�-�ĹHY=����ȍ��e��b�eŬ�Hc���}/dJ��4�R8碒A�3��@�y�i�9�ȱ�Vq��th���V�i%C=��I_�c*-�%��h& #E\�B��eӕS�=�N�\�z,^��n��@ Ǳ�C��w�_�
f|!�? /	�*�V��L_����3�L_cX //��F)Ap�k�w�Qy�������"���Tc�*�m�[��Tk�fN4	@�.��S߉&����Z��\��W�$���k+�ez"�����«|Z/?-1�伾��L�t0�~�9�"J�PW^���9^a���A&�����b`�Y���-]�$@z�,k��+V �ߩ�������r	�B	C��H��h�Q����,LZ`#��f�n����df�l�\��!f�6TA�D&Q�!R���1/���l�G����}�[��cf$���I��u��6|���ܐ�l(��VHQ��d�96��'���N���,Zc��߽�-�m�&	����^&~�c�k)kM�{1��_w=ڪ����]4CH���o��䦛z��S����/uz0����Qg��QS�.����hm��|;�t0��2穅�k5+�1���e�#�&���8�4L����ϛ���[7ج�r?�g^�_�_�K�w�	�%>�$��3���:�`4BOd#�)�����n��`��b���8��$��zQ�eɼ)/"���&_J�ʶ-��1��<�AT�8�I>M�('SUR`�����gB=��2��ږm�<�:"+/UOߏf��	k�:�P�z&�>��k��{��7c��'|8K�b�����c�H�-P 6]J�j�6��9WGyЦ��E�z ��L���$(�R1^�d,?��Ԯ�j�b�SC'���y�}t]o�>��N:���cW����T�zJpXe �vn�g+QE@-2�̺��w�� */v|�ï]�H2��MO\�/嵲u9*>Zl؛)��qb���ZC) �H�䗨�VwZ��H�;�ecY�gff��|��P����<.��YPL_ ��~��[���I䥩<��g
�g(�����ڐWA��RXd�B�倿3�V_Xn�Z
��d�3翇M}d>x>ԇ�H�>xfcd�����A�f�ս�����J&�?l���6��w�;8�^��hљ���<��*�Y�q:Xd��~V~�1%�n�/�<��ߗrO˹��4�}0lkt� �P��o���O>�˘1��8+�p����S�i[Q��	��,���X!���ɭ�5�z$ SR^�."x���P��x�hJ�Ѻ�O"��:���0Y=׍3��{�i_ظN�w��Bz߾-�ŏ�����wT��}�e�yr�E!�tM��bV2@{�q���_�r`���h�k{Q�D:��Z���^ͣk�K�h�L_]A/B������X���f�ˎԈ�*2w�?�2����}�:ٳ�`�(p�������Ĳ}�~ʀթ��JN�:a� �E}Ca��.$�ii9H&�D�V��7�C���Rh�=��W��Tվ�3�#3:��A;>=�ϠowD�@�	X �;&�N�����v?W9�ʔ����3}HŮ�W �報�cf�'��@^QW2�sE*�YON�[o�FG������A�p�-Մ��{*�!H�a/�I����[m��2�wBE}�-�1�8�o�}P�{I/�	�����zy���]����+�ở��L�Ң�'�n��؅<�1��N�X��@��8�-p��R�1@�A�SI|H�'�@���g�N�Dht�`�:�,�\f���E���.^�EiX�dظ�k�j��QJ"?���6D��(V	�H�c�A�{��X�+��e�a���{��M�Y�J��Y��A��Q�iz@��҄��f�f����d���kG��5*�8
�y��_����_��Q���]��f;)�{\���2��3����gN�~R0��*���Q!��*~��R���*NHy�Q�_V5|�Q����a Z����4ŎZ���B]���;�4
���)"o�=Aj��V�f �Y����I��y���h-�/��Sf[G0NM5�ӵk<�#\�����\���%���[< }�j@�Ř<pgx��*v�&���2Rw��)(�@� ���χ^X,i=_I��U�
7GM���m��,�öo��)�"1�صC�.�6�X�\���3�H�A�4%�|=�$��A�$إ~7�lw�6�\%�Y�G�^i۩o��r7�,*(��b�݌����p���{@�^��h���ưų���'�0٨�5 5���%�}La]��$R�I����c5^!�\��_�/�-��	΁hhʯ¤	@z���<�]VZH��8���(Z�[Ô�UJ@�Κ&�A�� цv����t��s���6���\q]�Xb��F�VGEO�⽠���P�~U�wP���Q"j7��^�e�[5���/ja�x;U����F۸�o�b3.���<5�ѹ�L�{H��齛ș� �O%�A����$D����
[y|gE�Xu���Y�G]׵t���63� u��s����$�2HL۔��6�C�0T��a)+�n����/,��G�a<�YR�!�ԁ�	��Y6sΠ[��z���5 �V��B�L%!�uH;.�I�BS�=5��rT��zL������԰�ȡ��M���#-t`<��;���!�����'�� ����'��ƄxG�l9g��o����N��x|�I\yٔݖ��@�o2���;a� "���}q���^%7�����><�F�AK!<ݱ[֘� �{�