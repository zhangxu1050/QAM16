��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv ��i��X��s�-�Q?F�`Y�������� I֏�׋������H[��9����ۍ: ؕ��6ж���Q��" ��y&���Y	6_���.���M�ݟ����k����
۷j	���`a�s�Yot1H���\��5	���1���d=�� ��l5�yFk��Ԕ����c����]t�VI�X�-;�V�x��৘:�~��Х��ִ�r�c��F�JV�f��j��/�����=vX��a�O�W���3�g�eK���5;v}aY�R�$���k���u�m��!��@] .�^d��0d,����N�H��7ǌ.��]��V4�񏣺��!����u��>�Mw v},e���yHD�з�K| (� �<®_��8)�c~�!����sW#-�7�iɛZI�D?�
�
�R2�;�zI"o�m���3 {y�%��f
�0? H(�몇T���i+�j���#w��P�>�acf�G���ߙ!\T+d��P��e�V�_*ͅv��ٞ*�@���A�,C�
�>��(KYr�Uĕ�¦Ec������@���� ܻ�aQ@s�����������i_����1�i��cv�x�o�ŰH��9�����x?�����Tb�ʎ6����l�k�V2
�-�O)�������Y�,���fo�
6�ś�?���u'_�z�cA��#�x�	,��X4�(�ˁe/���:L;�H��>H���Q�M�=7-��N���H|�lK�8�@�w�x�Xz��>�c	�����-�h�_U���G=t���Fc��5��JgBij�� y>���p�e��jH񫪁PP����dƩ��������=/l�=��$�f>@�Z8�%Qe�I޿���4��L0v�g:b�KY����C�jҒ�Z���%�T��Hm3t�L~`S������$�lS��/ �dC��P	ƀ��*쒻���"�D@&��<O����I���QY�¼?�������q�8r�!wL�S�AF�T�B� �����+N�K�ՏRЖ	ɬ�tn��I��N*X^h���S�&4h@�5�.��Y9¬����c�����]%) +������̎�re��t�7]��|���W,���ޥ�JU�)M#���\�s���}"^�Z�7�$��	��YՄx��G���sf�7{���A�Rm���MU6A8��EOf��ʖ��(`@5����{|�T��ך����񡵪x�����ƿ��>\��g�Zqw�c���rڠyHC��8��>�/3�/���*g��6�^�֏!�+e_N�����X�
���	H����@GnC�y�n��~���z���	/�~Į}1+���%�U�e�]P[ܪΠj���#�Վ��;{�)2��<ϟ`�x�)���K�ZO�՘`:5�C��;�$��Lv��^�	�>2P١�yM��&���R���7Pfj�A(ڱ�#����η]�.Dج�mDK��E#��KOf OT\Z�e�a�0��!�a3�&K���]����hဨ^ȥ~�51�	��.����$��dk�A�#Csda�"(�~c��*	�Vs����fz�����7n��}�@G�)����KlP?�x�G�CdC&g��.��P��j�j���O��ɇ�3�m~�ׄ�r��˸�8q.poc��L�}��Ϊ�5m��P���c�*J�*HP��tx W����<�u��Ր�C:�h�C�f!k��wR���q}�K�F����hq�<����)خx�0o.qҏV��+�e��4��	(�*#D%�G������!ig@�-�Q~�Tq��;��oP��M.wX��R}�������M#A�`�4%}��vE}3�Z�*<��_�<�����E0�W���J�œ��ة0q3�1����k���$�܅�CCqzn�?-[!��h��)�b#�h��zG��*JHJ���-���Y�0��g�YJ�M��6 60�[����⺈,��E�*�5}=�!^�_j~��хFD�^.�̓ԦT�
�o���g��F�iB�o���n����a��>��B�OGۺ�3�~aa�%ʦ���Q,�Ъ�ϴ��R��h�Sa��߽Ձ~�;K��4�l�Vy;���[�)��;���f��&�^G:P�F�5�%�7���8R��>�k_u��	 6�2 �}i���n��7�^^Y�oV+侗sbVd�h4���HX ��u͉1"�d޼-�{����`��@���V(y�~U�S.��_&��4�(��T��Z�\�{U��[�ʎ�N�ﺂ�$����Rc�;��ifcKхntc���܋	��ã����@��"�)��qp��H8g<�M��I��u�N�"���>PuL�JB}�2��`gk��ӌ$>��e�%�����U��
��E��% �Pm;08������]�PN����8n��V�����b�˫��T����f�}���ݗwm�YR��0���1�=���u��MSZ�Ůh�W�ш�:gX�'X�ɛ��C����(gC�+�>|LPH�8kN߸2,e�
�L������ajS�O���	�P��ۈdz���(o�iSR�.����s7��n��$�ɛ5i�E/w�2(/�UR���EGe\�X�z��b�K`�%θ-�;X��x�Pe@._*']����A�"xN��$#, ��/ABջ�%Ȟ����b�Bs�y�Xm�
ǄnS�gQ��$^4��{�K�]�����4�5.=F[�Ϊl3�E��7#: @-Q[iZ��q��o��R�ag�K�N�kc82��]����0�นq(r��;բ(c�v/gc�,k�㧒7�������8�d��r��̞���I�34�6��,�s,�٩_�v�_CUo��^��G�OK��B7 �r
��^;Z�%�Nӥ*�g]!j�g�b�i�2�O����~�p�-id�$����ΐN[`	����M����b6�����C�o5ܡ��J�ٮ^t�[���S�%�Y�Nsvm��]I�{���h<����C��y
�cA������@��M����*�~֢d���Y���.uD����lww�j�{��U�E�BB�nc��O�fkZ��p!�w��-��h?'��+�'�%�w�f�/�~ք�ȵNy�JlJѲ�z�Nf.�>��h�JD^z��E�u|��b3Yx�:�X�Kw	�>�󨯐�M�e�G���>���L��.�;�H�t�@�	b���i�]�������ٗ�X� 9fi��Q{�}Q Z�D��k�l�^���i�@q��I�����؟����!>t�K�{�o�D:����~�ؑf,].IcVф��ܙ�j�(Ҧ�T ����χ��ף����OT��%���T�?��ᐺ�4�[L�\��|͇qG�c�-m�5��cZ�_�g޿���\_7�G�j$f�Ђ�O���1y9e�eS��̲��e��}*Fy���L��~;��(�C���^;��:~���l�oe�6�^S����A4%�+k7x��ix�HYy[]�Q�Q�tQ��[A�8-��x ���)|��R5�F+�{߸ԙG��;DF���,�w�΢�P�&�J�N�M���*�o�n;g�Z�r��܋�
_����&�Nm��;�i��N��!}S��`O/Z���[�|H9��a�Ĺ���]+������B��g�����^KV6􁒙#�ܢ3�g�u=(���ܡ�!���P��JU���o����1btUx}�Z�*��V�~��@�)�$�� �����h�+�o�&�s�O�m�ֱ5�^�;���;2��R#M���P)��DTa����8��4 B �)���
x�E��*��ovBƎE�ޝQ�@����Kќ������'�YhV��`�ad�zb%{��Ӝ�N�S�T|�{���o-q
T�+c�'Y(n��	;��/N��M1�R�Gc#pj��!��2�x׫M_l�%&	���!3.���k;���؝3(�+R��2�󏲎<ARQ袿++5��/�`Y%)��?��F'\��ˋ�@���1��c+�yDrs��{T���%�2M��XV���p�V��� θ�0r������A�I�@���M�؎�lZ����<P�	�KK�o���/pvz�� �cxp���?���.pҳ���i�s[
R �@T)MeC �I�	E@��E:cf�-���F�� ��p�f�e�X7p�"��
K&��6?�E	'>,g���hX�T�3�1'�~^C�mh�N�&J�� /�;�U���|zs{:E$�����`��g �e� }�U�ǉ��mBZ���_�n�8��R�|Z�=J_K��m��^�s��l�)kZ��v��(��-�f0��Nxs��9@�K��ZXnj5�P(q~֩}L]���XGV�@��G�`��ӧ��!ԿHFq�&}�55o�(��n�tkD<���
���<�z&i>����P2ޭ�uR�o�x�H�Ώ[U��&�cN��"��� ��=�{9Z3cە�}���a���~�eb����8b���Z0��(���}_�v�Q��Amp���!�]*�	�a-_ޤ5��l`w��;��Z赯��u�Y�Q0�%���R���Q�$Ъ��Wj���`����
ͺ�A�4��{u�U	�>;��{6��9l����������?�(���F�ˬH� ż���||1�,(��v��}��<���$p�O�OC��K��N�DlI1 �3��n8�;
���:js.v�>����6�MIF\��G��(����~�p��2�eQ]`8āg�µF�& �x?���5�f��Ќe=���X��ݶM��1�8Jj�J���~I�/糡Ś������[����%`O�"�n3��uḯ���gTpcz���Ȗ^��`�0�Z��4�
����hHطAN/�S��_�����Jܦ�Ť�&�X�kg�z��,.�/�S�O٦��56��u�
��Eno9O�ؗ���?9|�M��K�gh�QIY�����tU���Ml�lWh$���5�p�/�:`� �t%�O��@B�����owY=TدX�)�;ʉx�Y�L�����z�r^=�j�ȶ3�*�i�;���R�鶄��[�Y!�)3��,��]�إ�bH�ԛ(}d|tY�����6	ڻ��3z|7`��Ԉ�IͲ 4H)2k�1���y������) =x�'Q���N`�(�<2X�-s��8{PaX!�]��w`M��ǎ��mX��H��U�MC�c8�9�=��ۮg�|��7�jLj�����+�R����J<����O��Q�֕ӡNN�����5�cd3]O=t�=�1k�uU{~5�6�m�|ۺT%�$<�B��;ӻ���9��L04-�a�i�E�Y��^�/��j�Gр�v�1!���q�	��i�1�-ߟ_{+�3�s�5U�B �j}�`aC1�:��3���E�:@߁�}�=�-�B�h�6�vt��Ç �s����OAu�E�G0����H/��"�[�YR�f>(�Ѫ�*�G����Bl7�EK��oT����8�f�iUg��K}�ɖL8��H��?�{�3����>.���VŇv�[�K��p��y�ư�pf��WL�+���/`��&M�ɚ7wDW�u>��Wu�qyB��ߎ��˩��ru�Bg��*�En��IL����$��ߔ����=+��ƩOgr1`w�W��ڊ�`δ	F ���
�<� �ިP�h~���=��ou��&j��*�>�.�Qޤ�fw\�f���Λ�A��4r~*��n�v/O�Xb���=�"��\�ĩ`�[LA)Rdaƃ���+j�gR"oɡD�E�EAo񩑡�~��,�^�4��rF�:�q��%\��0�kRi87��hZw^}J5'!8�t�f;Ӳ�s���I24�$��Ǿp��f[�C�k�}	�0P�	�tc3>@����s�yp�n��
VGt���*�
�L*weIs�~�x-�묬����Ov>[v�?�&/�ӐZB3��`}D����p<�o��Æ�;����HWŚ����a��E���4�%6"}\�N`C�84�O]����Ԣ���u��o;v-��4ߎ{d����4Y@��ɭ�Q�CR�Y�+�C
���8�>���ܐ.f�P�5��j,y�����hU�����Z/��gH��W���ab��c%}�Q��ߌ����f���B�����G�M�$�#/�0�^!�_�6�X�˷�_��BH1Ж�O�ysa�d���nՙ/͠��U۫�.�@��u�[�[����o`�?a!6O�N�ӣ%{���O�3�`�b�%#�CF5X�ċ�Q� fq%�%L7��ͽ+�ƭ�F��݀�u#��	��1��@=��ݚ�9
��b�S��XO�csQ{s�!�
Ђ.mm6�]���;�;\�׮O[n`aus��j�[��-w�NȲ+��)�0�Q��@6"ն�x���Q�?ɻ_"�M�9�4N$u[��I��S�9�<@8���B��h�`.��IZ�#��óKA�7F�~��X_�HQ�0�lT�iy����!8<U�
-u$g�}��s���*L)�yT�|�L�~� ��.%"� ;�4	��J������3%���g_k�]�KU��N�h#��~ͼ<@�.�PX�j�Z��Ϝ]6s0�el�1��� �Z������B-%_���j�[�
ֹz��\��hl���;oM�Y��?����u~́��^�4�#v���ր%�0����?e�rI�V������蔈%�e�Zd��P�
6�6�İ�
ۚ��$R����	G�Ӹ�๷{��2�A����ϫl�@�����|��f^s{�Rc/_e׀��!�TYDY�[��n�h���5M��X:�I�H��v��Ț�*GhE{�J ����8sխ!��9w(Ԑ.��i�#7J��5&��)��E&#��掝ѹ������'`�B�w)>9�ɋ��*�g*����NF�ʆS\Q�U��R�z�
».YV�s:�u K+�	�7x�bJ��J�I՛���X����0�~��pv>���tv��E��R�H��U��O�� ��%���9L^�E�t�٥G����lmM�ٶ����+ȴ/�-�����[c	�W',��gak�gX��?��sj�&jb}����� ?9�F�{��M3I���~z&�`����œ�>�??�l�\{�&��[}���O.Lzt���4BlIx_iJw`/����#��`��<��>�D�>�|HZs�������m�n\S{�	&���f�O�w���ZƂ�9@OQ@��8�'����ep]�R�1|%A��4����PYE۲&���78�vx-�dG<�5�i�t>5�|��*z3�rA\���~"�y���Y�1p(��'L0�&�Wr&��+�L���^=[��g3�䋃��p���� �s&V#R�.���ø�%��B�ś�K>R7� �����~&�(��<�#��F���?�J�0�>�ʐ��|Q������t�{��g&���Y�*k�Ĳ��Q��0_vb��+J|X�>�[	�����F�a���]�g\!���
1���1��N�.巭��u�E�I�����%
>�l2�6U�~���xxr
�W��c�S��O�N���ߨn�Œ�p8�qkd��k��yPR ���"s��xϮ�F�C�v.��Yv���4���>�L��Q`[&�׷IU	�^Hӿv�Wt�`�c���
	>��.�A ��zb���Au!�Ň����Q�L>l��Ly�Z'�SO����tVa�_KC����bm>��, ���1�P���D�엳>�f6�U�x�qH�5�@�c���&�86	������Z����c҅,����r��E�G�s5uW�G�(S��l_ �Y4��E��YY�ɤ�1�s/ꦗN�A@c]���9RU D�^@���n,�>�,����°���3)E�[f�;d6���L����ӏB�z�[��0B�R#7�m�"�"��o7���m�$ 6�6PF���/�܃)(�>����
k��%↚�n����QP�s��O}t!3@���0?./�	v���?M�w݇��u�z1#靘�[*���OPXq���I��9c�
�5B���E���>ί.L��E����~�ݯ��%v#��kd��.|MIUkK�uJ=cM�j)��]1G��ծ���t@��B��g�cK~b.�k�אQ���s�a�:󎽧juB�/ѧ2i�e��(aG��As�:���W��r��]X��sVY�8%*䠜�z*�y5S��K<+B�p������vnp6��]�(׾�F��V2������in �J5���{�)�Zi�]e�B�g�O�1���z�Sؚ4���JT���*�q�R�J�/�Q#W�{��*���sQ��Ej��C��p��t�Nw��v|�cū�1������2�cc����H���q3���/i݈>o�.��O:B�@!Zf�����Xc�����[�_+��ڥb6�	{P��ok�����X���=�5ګ�����}]�w���т��#�@�/�����_��1.�2�吮m�Y�H�P��C�f�r�ʁ
�p�0bs`�Z����ebz?Z���qm�
�a���oڜu
k���O� m*?m6����yQ��[{yֻ�=�Z�a�. �̅γlS�
l�^��R YoHs�[UQZ��������}
֭wL�M�CT��0r	�\4��Ak�C:@T���^�n�6�}t���������?��Z.�Ρ�S*��ǘ^/$[7FwX��ɻ�J�/lc�2�4s
q��N>hV� ~�X ����:�ׂ��a�����/�B����;yq�Vd2��O����^��d*	�)��?㙭q�1G����<�/ĥr���z�u��v]��Ѧ�ä�.�
_����ưEVΑ� �w�E��� �z$�_�Y2 �S�,&�")�?��<m� ���H`�|�r(p����$��Į��D%i�L����yR����C�!կ({�M��hu�'���jS�L� G�@�4��Ö�}�ڸ�����hWk�I�"�=�	�Թ��m��m��=�2\�������6�:��(Q��b�˻_����w�O;2�)
=���_�B��$��������nԳ�����:b�M(੒��|�.+gb0��~�m�Ud��� ��9Ιw�r��@�p�_�$�("뚱r��f?@@�dT���qW� �(Ri6'�/�N�� �DƼ�Ȫ�g�A�[ �����B��-
5������F��Ұ��.r���
=���v��
�~��r~+��#9t#�cXˊ׶cckv�ڎ>\B'y��*�+�Mc"�P�MeR[�����9��PK� ��t=1Fb ��1a�-�"�k�!�ސ}wl4�!������/�K�7��9�6NR�jC�����jW�	�a\���ܴ�{e�ܥ;�����t�P�O�ٷ{oA�k��r,��Ak�<�POk�։�T-i�����"�<�W�(�*�l XSX�)��Mm����;�aϲJA��o���V.�w�_��XV�O��f��cP-�_4wvՋt�C�-��'��eP��:��i���:)�ת�Ip��d��■����),��.ʮ��d��u����ԑZ�êJL��{���L��x�)�C'�?��7%Ce��ߑ��+������m�	�H�Z�2]�0�/�� [�za�k8=z�7�m�d�Aq�u�bP)@S�q�c^9 &����x�g�l��.H}�P���s��凾��o��b�~z�[�+�;]�W0H��"��hvr���OHa��9���,�D(M�I˹a]��_e�= c�p5�)��oT� �}?p ���Ku΁)�4�l�@��Dg��l��afG��pQ���ዷ��ü��M�����S��4��a�M6���;�&��o�!�rZ��2���``*K-	V�� X�d��QcL��U�C�&R��{i�hTjZ�[71+>�R՞e���x�&e�t��b���Eͩ�/q�	<�������g��?�)�"��oj�K�G�Y��'��[���L��J��3r�*����ZƐ�Z�e�q�#�c�f�$u��	�)�H��ܳWN���@�@�a!��+�E"�"�:>�]x�6����#��"��춌�Y����&�� �0�>7�`���*w�9n�&H<�5y��o����[�~�a����SSNV!4e9�㜿�2�ɱV:ՙ�|e�O�
8Q�����D�c�wYNH&�Ӷ7/�����2�J�B�@c�CuLv��v�'<a���n�س-�$`k�����قґ�ҧ�c4�����R9�A���š��5Q>v!U��2�e,�%.����Uk�O�OƆNł&��6�d��U��JcԤtoC��� 1ڻ�*��e���SD���)��N�R,����CC�/���sGDO�e�O��5ۙ�G��iI��,�Ņ1.\��{��]/�@t�1��i��Z�D��7���k��{��9��Ŭ[?�"���Q��U�L��c��I��G1�q=����7�U��4~3��*��؈��\`��}���֗H{(y__A���Wf��H��~8X3~X ��r٥�ت�ddqu�����	�&3RLl���z)��_�Y��k_5O$Z�@���\#��t�?�yg�>����7�X��uԈRq`_H�h$�oH+�&�g�EؖnMfn7_�l	u��"��F���w��/r�"���:�iR#=����P�]U߷��ruM���� �ԏ��^[�Ղ����\9P�W�ܰcIA�H��ld��>a��X�w�7I2�D���x��@���s# |������]��c������+|�܀(��A��Lk
���Qd^���ѭ9�S����:���o�Mq�0q~�2:�}�EVf&^ ������Y�ߏۅo��Z��������k��҆_�;����3��I����l�8f��M� +h�߃
��X7���K�{���X�>�Y���f��/t�xS�����p?%T�� X�n�vr�N6��J��3"|�:-w�S�g��0B�=n��h~��3|ɾ��;�%�l��� ��ɼܾ��%$/yX���qSwi�u![[�y�%��k�"��w��_!Jȇ��<�:u}0v����U>��'D��'�A#{�=���cQ��@Q4��ar"&LA���ZAW���GyY
_�Iv �1ˆ#���1;�ک��8�����ʷ�;��^f�H'�T?��;�C�5��;O���i%���T8:����9�g=i<�׺�@g�A��#2�B���#'�������+��2�=\�O8}?�Kw+��,j_��3� ֖A�f��{zj!��>_�]0�X������0bP���lFK�4��;��V��٨��Xa�E$�>~�7B��v�eh�$@�	���!�j�%�z�'��B�d~�*y�ߖfO_`, (F(Ґ\��z�ʑ8./�c]�]\�������gO�jjm����1����D�j/(�a&�nb�B��_y��W$�.��� F���t=��+��5�MĳTA��� τ*�WL%��B����@��Kq#�9�eC�X�ʋ�q����dX������M��1t���o��}�2�r�T���߯�"-^z���"�Y��5���ss�u���4��io����J��I4�{���X�H+��h��9�h�%��)���Os�rm���c���U�͎�d�v��V�㓌뫧&��e��xaR;V������)�%�[q��i���]̣��6�ϭ݁W�Ҿ|��k�,�/Pj���O��.[/ss�`�`ccbT�f�-��1��z�"5�3�[To�� �� _O��k&vll�nЧ�(�YG��L�	1	S��!��k�jA�Г()�`���v��d�ѫ=��3A!�o�-0����<k�E�l$��l�gҳNM���I�	�\ހ�b������P��]՞��aH�^31h�mr\��l{�)�m3�$*�����wK�L�x��c����E����rc�+ů_`d�.�̯1�d�J�9]U�,}�(q]4�3�O����t2���<�p���ݚ��}��2"�Ǥ#�nq���JI�!u�[ؕ��/K����S� �X�5W,�S�	�lVÓ���0:4ں�	��*��j��]�؜��]�4n�pR>��6���=`k�5�g���(����jUZ�E2Ӽ������������$�����I^}��tJ�<:��#��P �`��hf"밁����&i��ə��Qr�--u��4;[PV
��Ј{�9d�?�-����)Qd�.��i��i~	T�;0����Ӕ��E�bG�p"-:�󈍹J���X�Rn����;Թ��;P]�z ȋ�s-&�%�t\#�z��07To���U(�$2TYh�gy�������b�,����|�?B�uo}b���d�ee�)ĸ���V@�hIh'y@/NS�$!@�#��j�DA��N-^�v�k��q.t_Zg��d�~�9�}~�G�g�A�HT�g�S�	���#��Hs�hN�g
�R}��WR�/[w9y:ŗ5���\�p�ؽ��̕�b�Ir����Ͽ$0�����>�@�.�UN&���X��+��>?�"N��k�9��x�ȥ%\�q\���V?7U�*K���O�Rf���y��n�[����;�F�
Ԡޟ��2��,��� �%��H�Цa�:%����v�U�-*Ft6�>�4ShDD��8�X�v����6��h8�S�L�����j��:�5�"،�-zF��`&�_������>��(K����5OY�,Qt@������O����hu4���%��|LJ�@E�vGC���?�3��%;���^�-�H�̫����c|O��c�� �}��`$�s�Q�c{f�
N\��&�d������[��]�`���NhB�����6�'��j��Я�n49d��d�����:"�ǽ�Eeq�Z��)��'"��)A3]-�5?�;�{*AZ�ce'����0�w�K��W�MW@�q�*|�i��E�Z����P^����V�j��g� �������1��_�v)���:뎛���p2Ղ��Q��h:����uX��W�$\�B��0E��QV:�������s�w9���mk�X%<7ؕ���R�q �h���,E�|�X#<š����<`�o�촙�ﳭ���.��}LD��Z�͎Y����%� � �Ӄ��9�.`�٬I�y�؄Kv�r�	'%��F7�x����^�l�`M�~���X�'��!]1�cwF��#�r���L�ooHuig�)[�([�Oj=���J�n�a]�KMc�p|}.(:z��R�j���h|  ����_�R���gY1å�M�����80����5�������ek�M�z�2�e\r��"[�3G��R��JI�E9����rt�+٘s�����L��E_ǿp6W��$IqІW��%	�~/�?2���]m0��Z%�	`�����C���Ą^��������N�S~���W�uDi�I�w���XF��z��dbp�殪7[=+�ִ�,Z*�\�?ɛ�"ft6%4=�� �,�5Z��R39�2"�RP�Z	ܕv$F`1tdeb�/^0S���|qK�P��W?Ƅe�3�s�G,X��+Ȧ� �`e��C���E�*�9�G;��Š�m1�w�ŉ�ߓ {P�?�d�����E���y�����=�g��(�f/Nά�;�孨����l����zo�(9{���g����/_�����6��xS{������Mv���vs����K�zPea�n�85�⽔��M?�/fX�=���;�]��*�rd4�G��.�S�a���|��,)��YA�<��� ����`�T�0���;Y+.�tF@Dw��[��얺c��1�M����Kh�*�^Vxn?�)�bY��Ϋ�&��Ӈ�V�~YѥF�KzP��X�,�1-s�B�"�b�����ҟ(��"�BݘPf�z=.O�W2*ހ	hP��}Ls�AVS�a�q� �(
�>�XKQy���m?9v]sTy��D����Ip�"�z��|�\���whV=�&�H沵;ҰbSg0Raܱ7��G�^B����i�\H����f�d\�m���\���Ja�o��C�-��(�Oc�9����=�ΐ�P|Z�p�<'�����d-�)�*":xp������
;�6�IX���Q�#���%v�4�p�'��U�' �/�h���٤ߗ�g����K�3��S�ڳf�y������͸�Jk	&�M�"��<DH�)�,��\c��|O�o�e�=��QP������~�h^`=!N�Y��C(vk�L�-�i�#sZY�:���U���߶k��bn���Q��m�Q�m1�7>�d�N�Tg+�ZU�vNat�����-��.`*K�:
XUnBd���Ҧސpا44�ɰB�{�3�_8����tA�sNy��A�x()��M����ɉ�`�Dr�B/����*R'u>Fl)�+�8'}� B�خ��1�?�<�b*q3��Y�=�q��$h~\��7�'nj]'~�%�c�I(d�x�������.n۠�X�q��\�n�a�f.��0(�!8�aw���!jT���R�*�-&�S�`�;WD88�w�kNR�[�秂Q�/��vg#-�RE���K�8���Tq�Jbu�kAk���v�,�{^"�e���0�# ��z�b�wW-_�����{�?��ze!�ë�������^�`�;G��_.�ԧs�Ue�_��H��
�81����!��0M��"4h�16�u� 	i@�b*3��ߪ"��wSN�J$bk���>�i5�s-?�|�+A����	�Xe�)����C��ӡ�`d��W^v���z��2�:��߻uB��1%�3|�i�)����z4T�2d���f���А&���Y�V�Xd��u�.a��F8tE�. ��(3JԤ�J�i�
�߻*"�u�/ �ÀΕTS->�.����^6��"b��HS��y_��H�Ǌ��C����4�`yH����;#��T%�>{�
q$l����]�����1�o�RT��Q�,A���];Ʋ̅a��.����vQ���f�J�)�6�ƸM2䨰>H�߰�ѭ���rǅ#^��]i��������q���<4p���##'��$�}W��n��Y�"Wi�6HS\���������.c����Љ�HmX�����/tp|���s���-����ɓ �X���7I����[i���}x�����j;��\(l��!Q�ERI}���N���
@� �Hy0���,'�dx	�޷��H�⎻_l��0��BI�z�g��Ru!��wH
g=rUm���Q��������t����ً[۳�!���j��T�y�Y_z%§~y.~���m~����d2��������A��?3"R�P�c�Ƣߟy����9�D-�ǲ��g�Ȭ�u��!�'���=� �Tȇ2iMF&���U��6������� �C:�w,w�p����f���*��p����������L�]���A+�
3�}��L�޴#�g8��%����fI��}���H�/����Y��7��b>�[�t�ⵤ�w�Z��vŲd�3����Eg)ǻ�7�@B�4%��c����x���SsG�0��/9��g�m�
A�S�w����d>rl�1�@��:�-��a��E�ν��}�1��|A�;�J�s����>��ق���=��)	t��e���R}o���'�.Nǘ���X��!�J,��3b�Y��:�?1�9[K������9�r�hj_p���;���'�p�hLuN��p�TOQ4ɛ�o�).�TuMtgIO�Cp�
z'5���2�WR9s��ܐ�� ��n�@�t>ӓ��)i+lu�����Y���{)o����=�{��u�v��k*�;��W����O�&�TO3�S
k�@`�T��'�]I�Ix��7b�|c���^�;�I&T#�=��^����w,�c�x�ܚ�A5J ���w!�'{� ��a���u�Sm=��Ul���>=7��_J�d~��i�!��ﭥ�����o�����AK> ��R;�X��SJ��LL@�=~�_�~�J����^`��3b�,��ޡ�
	��åj�,GO�	�E�\�t��9����у�|�����{�LN�Ìz�����*�%�i��p��&�@�pJΆ O ��S~�wcA�NQ}���61��u]��������=g������3��2���h���?�u�52<�/SR�7t>?�;;1��P9������Sy�W�Y�:�����Ψ~0�a)���yո �??�7���ؿ>�� �b�Ʋ���m�Tg��[��|�@�&�|sW�%<��U�1�㼓.qr�'u6� �A��>�H��8��^�Ƚ8�G�F8���z����N���7��x9�@w�e-=��a�i̹��^���	z�<�)�2j���Ds���]2~�_�Zﲧ�G�I
�G��J��P��B �U����*���h�h����,P��JԹ�p3�,��8%���z�����V�R@��b2~�H�8,�,���7�o�Z��H�bP���v�`�YK|���5)&����U�lEZ�
K݊����},�!""R��$e��_��MJ��w>w��@�%9?,�j�����k�Z8	w�P(8EN�r�ê=s'f�W��<��O�gb�HNU�,�W�[����pAI#�͗�uy�2�ހ�[o�\J£H֮�K���w/lɥ��
��eh��s�^;��0���x�C4��20֬�� ڄr,���o�\_�����3�Y;e��x'
Yۂ[=���X��}ÿ8SLyѝK��o�&&�|�K�{R��z��WrD��ۆ�t����:Y��z�9}��,��6����7��߸X������WTfgg�>�Nr��`g�j׏� ߶r��@�u.��l��J�L�$�G���\XK�����x#j�I�z^�VeSy�B�ȞL9���;���a�#�@�^�"1(G X���CI-��ur�n����=J�]K7O;�Ȇ�Xmk'~�?�+����Z.H儮ٴ"ǘP�R��-�]������|��X�M��HL�l���>[�Z���H��axկ���p<ir�39fL�>�1��� �Q礪Β��ڑ`�����Gpv�|{[HJ	�8�V���]S�:`D.�q��"��6��a��gJõ�?��n��| J
�]_��s�u2�8%w���ߙ��%�M�J<��xU���%79�6^�K8F��4���l� C��=���u	����x7�>��H�u̢o>��]�/#&��I�-���W�h0�%W��5Q��(�3��,�/����E�J�
��PF$y9lD�S�[��QE���9��#�_骏��M��i����i����+OU͸���R���M��������������|ؔ t��֭@6Gg�uӌ������E�+E�@01��R�|Ö�@��$���q�o�1��T�'��)��YL��my���X��!aK�,��PvO��p�L͸��Zȣki ī�sEV1�˶�O }gٱ�p>���;S3�lŇ��7�X��d{�����磹���y�Z*��&/��D�_?�&q�j��)l+DWer�ǐ�-�E�nP�6�Bu���%��EC�|3f���1,��rY��������=M��1[�ơgc��"7!��r�K#�tZA��6pe+]�Y88`�Kb\ry�~��4�����q9�Ј}H�xс>��A�_˿��
��9��O������Z�/��ׄ� 
F<Ϗ6���K�\̓�t�D+�����,����p�i��睲���F��v�f9m�<��(�����Z�ϡ5�#��`���wxR�^I�ok��:�Be�k\덷dp��	��#e�>���op�T@�!�b���4a.B����m��{O${�� ������o}�S&��z�^BO�����KC7�4x��=g4�C��+��)·���j����n&� A?I�u���흋+L�|5��R+�� ~߉���:�1��j�)�17>$���젰��f��F;Uy-~�^��T��ht?�G����8�Dl��u���_�Yەуl�����TϞאT�T8� e��b�O;w�)D])"�?�N1� ��m��Ŷ?c
�-����3q��A��-�Fݐ��Х�ָf�[2*�a$��prW7�^�{�qgZ�y�C ��'Q1'�3g�O���'�?��D��!��7�ªL|͖�EǙ��X��U��፪g|7��1;�j��]����w�V$[���������=n��{����� �x��ZPp��t���Y�f{��I�^k9�HxcX����-	=��n�b�^�zk�Ҍ���n��V�=�SI�9�8�Y����g^�~P�nS�����z�Y��O�sb�u 1^Y��v�G����i��z�L��Q�@�_ic]������G;�3fH�0�@b>�A�ӕ=�7��9:�_5����y�x�_%w6 !���f�к&8�1���DN�-cSr��R��y@�P�ר�e7�3��:���G�)'6�=�_��w���R�nh�����W��E�!Ggɯ!v��v�-�P/x�$J3e�d�+�R��)Gh>��(r!�'��.X���g��oa�l�lMU��C&u;d5�Tm�((npf����fv\
]��q����> �5<[dRS��~�*�-
�|���Ck|m�v�W�}.c&�-y�z!������H�s!��"]ݟc���v8���̓�˩�n&VJxh"���`��6;:���p���>c��ۣƁ�w�ŀ;�`���{�f�;u�7���**����F��p��V��a{+g$�)��R�g��=V���F���vL�o�d��27�����i�߫`�$}��#�좢g�*��Wl�[*m��Q!8���&u1�k{0�&N�"�E{Yd���U����|s��٘_U�� r��g# �1��i���� Qc�WIok)�A(��i�K�?ΞOv,$�7��1��+�<a�/��I����֕d�;D݅���[}#�l�H�L��-�5������m��~�7A�	�<��?��~/=T�A�^�}�~B���@��:3�8�g��16Z&�����3�@gH��eD{�����o�i��cȜ�:
 %��rw��ɮl��`>�n]�S��#���ݗA[����_q�9v+.�m}������[���uo�m�|�/�)���?�}Xg�5�F��2�Xg�=h1��f�?����]�g�|����G���6@�n�(ڼ\4�7B��t�bkCb@Y �>e+kp����ez��qp��弩d��$�,��=�1.���vY/��(�C��C������Y���k6Yx �c�c!�@lγ��^�iu���2a��hؠ�ˡWI;�="��5���H��L�DI��C���̠���t!#�}�x(j�ւuw=�����C�aN-U��TTe�$��ʋ��f^:��+B�f��9s� n�y^Ͽ.��Y�
�>'�p��>��RX�7 yZp�I
��z��)�ە�Mq���47��5�p�à���טӇj���B�l�����hm5k�25�,&r⧐Y�fI
8E��	��-�:�m*�a^!�I�b��_=x�Qz�ݝ��
	� B8?����	�W!7%Ω-4���G���0yQ�-3���Y�hҩ�g��˅m�H^�:��TH'� �oY#كL��A�C�Ɠ"0�i�� C�YE��`Y�8�P�vn�H8�P��a�Su�v۶���y�F]2�KY�'/�4e��K]�TI(���iB��w�W���M!��%q����*@�zf_JJt���}Y��+U�b�[�ƌ2�O�f��7ՠ��m3-���]s�!��H1��-��C���3'.��G�VA��a�#�ƹ���&�����+���ĺ�es6N!�zdnH��B�����&�נ�65�`�*�Ay��j֥o���w���F�ǙµF@莣�7�߇>R�����E|]�w�0��1��E[��uOI��Rn����w��#��������k����鐒�Mݧ��5�����r����w�0v�)O�\�e�5�}G��������k_F�h)��7���3��"y������I�C����da�h�;�IȵԼ�%*�f����N�pE��a���xZwz�.ț�ѓ[.���,y}:_����
�;(*�O���|I��7��ᜊ#�f���9e[�z0��B��E���D�֑IO�(&s�BG�7��CZ��P���L�|;�D�h�6�
�0;jq�ٷ?ݦsp��������0��}�u�l���j�Oz~�R�.���{�*���TLm�6)	�fB�Ũ\4�G�gI}��~Tb����.:�TI�݅\|]�[�2��H�cq髡 �+t ��ҽc����ЪV �
�*����-������}��Hd�E����jp�U�<�Hxo���,�����/��Ed��g�l�ah��ӗ	��+i��A��N�o�8��?�Gq�Y�V�ե,;� w����~�T���,�&4�3rÕf�(�b����$��א|�]@veI���U'�!Y2�7�#F�$ϫ�R��.����1��>mg��m�Ρ�����|�����9$��*�ό��(����Z�M���l�_�yu�y�kG�XL%<�~V�����)�4�54�X�9ES����b���,���2S�kpU�;|pOn\��F��Q;N����:|BT�G�TB��I��=n�o(���X�{$j�T�N�^���G��{���{�6�nG��v�;��=Sy(�DS��?�^2!e��M�՘���9���.$��z�G	������p˚���v�K�`<o^EqqO��q�O��4i�w��yp�
�����;���6Yq;ֶ��p���C&��� �Pv��΁թTr7ܐQ��0�C�Kvuq�n��g�I�Ί�{f���5���.�:-��A��4s傧�$6"��qU2c?�>h���T�Z6z;R2Ԟ�j?<�R��i��Bxy7�}.���g2��-�὎���<�3 ���B�/N�.w1+�^��(��gХI�%MD��!�%����k)|Ĥ�"�׻A�ьw�o���f��j�3�5B����P��z��	�{Js?3�����?[���\m���PT>�eց���EG�7'�hH֗F��N���z#�g��:? iJy�;�pö6�PK�8L�������RԂ�����`�j��j|mV��*t��rCT}ը4�Ya �!'�;����u�|���b�O8,xt�.��8{�qRg��]��]{P���U�'��7�λj��U���]#r�����wnr��d�`���ܯd�1�>��B+����D�*<~	�N���Ӫ�����S�6"^�F#0宕�be�z��п��,6����S{���N�4�����g-�vW�g�c����4m�;�6$-x>gO�G�x�P<�M�k���=�8�[`�^/AV�~Rn��?ůy[*)1%W���D�\��.���m�HX��l@�j������L-���yȝ���P�����'>!�ZW"�Yvi2Y.�Iz�ԭ���؇��i��MZ�t>hS+�nRX�z��ϰ���JvYpʕU!����Q�&9�5�P���,�@2���]�,���+0j=$)nݽP�+,����p�5�.T���4fg�?8Z=��ĔFXk�p�^�-c���h۴����˄Ȁ��*i\�$BK:�)*�[-54ym������n9)F�s���N���M���%�X�q2h�U
se!	s���Z�����&IWC�*�3_����h��9L�'�;�[Y=*��T����T����q������?HG�P�<2�)��g��z�|�?�=�:|�e6��Zj�
��UC���f�e�6�o�K=ٞ}C�ll�?Aia��w�Yoɘ���v0��p݅�B��r)�����;�#�<��I�~��|8��l���JVK�-KY�f�k�Z��g��j��)�Q�J0��u�=��X���M�G�-|2�-';y��b
;�aO�,K� 
�V)�M8�����_�VG�-���^����R��N�)j1�"O��{��'���4Ց��a�_��DN�ul����Iģ��öE��z������vL��6��<�M4~(n6�TՅ|��Ƚ2��zfx�