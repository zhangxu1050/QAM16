��/  �-yfJ-
y��ѯ�U[�����V_� ���rq���~����Į����s�A�i�Q�#׏���ƚ���}�%�ǌ����3ؾz{�C+*Q`I�l��5@4��m��ș�nA��z��xc1��^wY�Z�Ւuk�Z�`�x-��3=~9I#��h��je�t{&�-�O莜fF��J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&������*��q5Ji�6�A�+�Ak�ŗ��Z�h_��f	}�G�@����Ԟ�������f
��kRN�������pm�bGCA:T������Z��ޗ9�Kl�
�f�ⴷ�����s�`�@����X4( ^v�UWP;���;75�U�
�\g�vC�HDM�&����H�i'�������>�M����n2fч$42>레Xɲ{�7�86޽��/
F�eQ.�~��O�rꢓg���@���!���@�:m?-T�{/����=�y7j!��#)_��A,gS{�G��,�1qo5աfK�b���БOJy4��&���\�Mǂ�zH��l>�`�J�.*�@SA��-��p���>��]ήq��,@�5vzV�����751����3���]��o��ڇ�P��D�d��l��t�3I"X�u,N"Z3���ҽ��N�¦g#I�EAR�>�!�O�cl{:�Р�Wtx��5�$�9���&Ha��(�F�ajk�#�:���c�,��f�A��,m�6�F�]%ү��M.0�%[Q~��A@y1=�����3p?��:
ʆS>W�wC>�vD�J`o�h�������|20t�˥����8G�{m+���m����R�M�:�葋�W� �E4�c�>���K���nHY���'��?Vщ�"p/�ysm�;7���l��
���&�W\T���y�E��w�S�>#��G�R�A�)i����5��CsP�0/�)��M�ּBO�D+]MW~V<��h�7/qZ^DqB���_��?��t�5��;��G���:�y����9)����������!b��ّ~]r"�j6���aA6�T�����R�8.����O)�Ļ��0���-TE��I�l��T�<��Ʀ(�G�&��	��L"�R�J�1���S��<�YrZ�K�q�l8�8TJ�e}�EbLZ�?M�[���j����92�rd�͏�n��z&Br��mV3���g��=��@�𦈇$^_'�8��e!4�g*��Z��8�5�KܢYJ�o����&��+[\=n���g��1u�0��=�1M͓FC�R�qz9Ƣ�)��i5诵���}|���C�J��CTWl#kFM��潋te�
_Y��!U%����Ğ�go�J�1�ңx�o��&jĽx!�������ɮ;f�:�M�tFF�I�?�\˜'�ɥɠ����;��ᶉ\9:�9��&U�y�W<�7���g�}}u����y�[h=b�-Tɍ�ND��kVg�7�@Jm��
�lk��C�4�8ÛVntY���yk���i� �)w�Ó����2��t�%Յ@��s�B/�/��G(��(I/�C� /���D$��o�S���
'�Oy��,*Hy{��і?�;,��h�����ͤ�O�z$��yqa;��}�|]��4*��X?#�]�%��o'��e�F�f����}��� �˞���N�G��{vOdf"Qe��w%��,�-�"t���-�e��9ä��wa-c�Sy2JQ�
�:e�n����Rx�#���qڧ��\��?Q4^��W��QZVq߭�O�G�?ᨨ��DAhcA��|j����^�:��X�B��(JY���Wn�-y/L���k��)������ϥE���~����`���T"�FJ9� c��1
�pI0!�.�|ZXeޔ �"� ��.!�m`�Q�Y�{Ri�?��^��>�T�[�����U��T8|�Tfd�Od1�$@�Q}��Mޅ�82�{�9�\��Q}��o0��-<J��	�ǌD�&I��q�9Q�c�1y\�#|�k�����E!�MI�����k4�B�iT^��|�j��9#��ZF��ᨤ�79��
��f��L��iV���k�o����x{�D�򭈈��Vv��K����N�	u�K��g���m�`>��6��>צ{��m�O�2�ڙuH[_
�]�0���]&��}֜��nl�y�b��T�_�dn����Uj�"P������-�eQ>�*�����S�k�r>4kO���~���l�Ҕ�p�@U�5�vk�ń�9�4�:)�N%h�?�_�����f��Cg��K�s8�o���?��?��nv���Ըd?�#ɗ,��������Y���n�� 0~���&�D��ڡ��4���x�Ǉ��̏�Z8�`�9���c��^�W%F�,��=���k����e��Y"uI�[Y��;��#�#�$xA�`�.�I��	7�X��l�'}�g'xVU�N�"���)}�5{���%��`6��ʴi�S'Q�~_�����Ը�,8F����U�q�,0��+��e��j��Cڤ+�9G+u�����c�U`<�����OSF���+�$O�߼��$u���U�̲���H�����~�� �C��q��D����MG�t��]})��X���U� �����?��V�e񨍻H$����xx�葊�b� ֝�EJE;u1�:���wK�K�']9x+�MDn-�wp�C?�TH���t���0R9�@{wAF�=�d��lnFA���>��H���$��g�@F�gu�c(=��Y5CkӼ"��##<�avjd��|~�y�9�Ktm��p����a�֭��}wnW�kFD�lI,Y��!���Cm(�%c�z�_[(���
���	L��H�f�B=�!n~�٬���u1y��>�Ф�Ŝ+�����]Gz���Y�~��;�"�9�B�kI��C಩.����Z�7�z��:��VR����iV���m�#�r?G�VI��4`�R�u%��1þ�\/t�8���F�2�`W�J5��f�V�J�4�ՖP������h�0W�P|��;��/6��c�І)��&T��$����dK�D�n�6i=xc����T�,{��D�	3�Gac���:)�d���&oz��gg3�-iۙ�iNJ�W���l���F��G���(�����f�*���R���P����n*�b���_%%b��
4*o��s��S�wwޑ��h�r�N,mqj��7ވT{�J�`�����Ǖ�t@>��`hr�I��E8��]�N���bch�D��e��[�.+%v�̵Bϐn��]wP�C�OMuO�H>�
s��Np�!KB؝d����Zr�2䘔NſA�L��wM��������T^P�ʃs�������ދ��V��,���4���F"��G
�P�q7������\��:ۚ2�����	��K�;���һ�z�Ŷ�I¨��+���x��_�[�I��Dk���uJJ W�x�=�6��JP�u��m���9y��A������^O��2���/*7ĥ���yS���X��2�ܫ�wm��Ǳ��=whrִ���4xM���<�=�1K!�P��=��d�1��j�$�?ص����R̻�rL��Z/gSš�s��n��f���Uehs�΁ ؁�{�bO�4�!�d)�#dOl�̧@�o|��آ[Y�`��^Q�����dN9���7 ՚���yh�`��H&�,qe�z
��9"������@;��?���P�lu>ڧ�1'�e@ݻ��~�n����TO�YT{a���\;mF�ۆ)ܷV(ee���uY�.��G&��N�m��|Ȁ�B�����PJ�Zԋa������j����m^%�d唘=��<	�ƣc�Psq2G�~��>��>�Cu�[k`�LU�4��k�ɼ4M��3g����9L�.��S�����8z,������
͙$�%�����2O�~̆��H��9w��yk����X��*>۝{D�Tw���!�/�}�1�U4������e�`�*�6�y��+��-ٔ	i�u�����B`����$�����أB�������H�Bi:u����ú�V����u`�U�){
��tt��x�t�K��^�Dҝ��\{ ���f��|t��lJ/��d �7��r�mO�҉���A�O9�l��T�����t����HEJ�ji��#��v���#�V�a�K`�[�S�+�l���ċ,�8�|J���>��N�9.��EA�z�9��;��؍zF�IV19j��1�@b#�e��- �VA��w����*�ϠU	Y����� ^�V�Uµ�%&(W��S�ʋ��E�����m���F��_JՖ<�e��0g1�w�x��[c��]&D����|z'�;�� 9Ψ&�<�f6�s���KUꬁ��mR�ߩ\�3�t��^2|ZfwC�s����a�ȕD5�����47׸w5$�O��[K��y��
,�S�9RS�h\��k�P���n�Rr�����N��������)�wagc�i\��?g���%�|��fQ�w�"M�0j�HyZ�biɎz��ϱ"��'��7��4�H]�(*}qˏ��x
KK�i�M�F�`>�g���5����,p@��Kh�{�d�HX�x����)*Ŀqw~?�Β(�˷m�dG,{t�U,p����T]�0摆::WJ���SN������O��~���"��On�aZL�����G���G�6&�/�>z��� �hy ,��9�� *׮�]�,y�)+6l'��HK$�V��}���_����h�����r1���6't&D��<"�c��y
��c�q��C�7����~@y�J�|��t>Kh/g�ƌ�ocתo���(qc��T.3FNy�k��h�ms�iF��#A�����l�s�\��ֱA�������t_?������w�Lw� ��YֽL[����n8H�Zkl ���L�d�}�&���Үe�/N}���� �����g�PX`����tH!H��_�g���E�\�x9�`W�9£���TBX�W̯���"��`�����Tc�"�U�Y�,���d|qٖ �n#H�ˇ�s!�� �Q꫚�Kwhj�Y �eZ���z�P&�|9���'�-��I��һ��>Kv�����xxod�]�_��@�d&���\.�����d$=�NH׺�����G�a��}>�0��+��]��tx�5J�帺�p8>K:�_�`�X	���r|kU��O��rq�� @.��\����sWV�N����h�UG�SM2�M[�1�y� �A#R$��M��~;`���_]]x��	�W|DKӇ`�0�"�L�����FJ	JTGS7����䃑��%��K�a�Z�.O�O�k*ouk��'Mʺd�rO!��5 �%�������Vu���S8����Z�Q�:O�(;�S[��6�Umi4��C�]��ä��&]�*�%��'Կ�yC>�:n{�����xS����`�C��GV:�"�_�6��Y5=����u�r����m�l�������h� ����fW�*�Ok�R�fv1�� �8[Y�kе(^�'p���.�:Վ�����NƁ�ct��`Hώ)�fO�9	�JZ!B������d�|;!ꟃb��:#8p'�ƏK��Z�2�Qo�{���j#<����;��k!�6]Ī���3;��Yr3�,k����}�Z�� ����b��?nҫ��K"~�={F�NU���I�:p����C���2G�B0������}Je�g�K���΋^�S֯��������r�%�Ǩ���o��Gj�������*�|49���\ ]6�,~��|K��w�:���
кL�W�n�!���>CI?Ȉbt��;(���R��������d�){����Vxs���r�|��f$�#�t�y��T��	�����J�
�A�rZ��;��#�u����v��\��&.�7]E�Q��o,9�-�'=�n_AU����Fb6����~��rq�ͮ!̚#'�1�����bh(Б�q�
�������[�zZX@E/�������S���'m���	-/Ś�H�=�gM��..U���(�aI"�Z��D���a�9(�ܜդ< Ce��9�W@�)ǲ��4�^�O�異kE�΁�YNՈ%;�g�-�R�IM������Q�"o{�]_���gK�bG����
K��X�R�[F���P���qi���>�B�9�Ѳ�#����F������1;jSSĞ��$!�����?U�	��q�:�k������{c��"\Y��	� ���J9G����审��	ا�������l<(���40uqz�'�U�x�C"J���z�vA�}e|�m~*�����<N  '|h.ێz�������Y�m���A�뷪Nvt8��<����w�lU`��[�xۄ(��w�|��^K�녏���ڪi��	Qv1iܚ�U-�H��}�q�@�bTbM�e,<���:pa5����B4�Y��Â�Wԍ�$��N��yIR��!6oy������^��Ƭ�!G�Si���h���82y>���S^њ����MN�7E)��ˬs~�$��Ⳗ��)Y$��I���0����qvz�C�V��9�%;�R�%��.�H?E�3�S���Ԛ�7���4�����KK;�����'��y4g_�t�=�R�`kY��V�;	�/Q;���HQ�Βg��Z/�@~�a�|𔨦��=���O�n3(M4��/�:�P1BU��2�V{6u�p+�$l}����E)��3]?%�I<�D��(�֞y69�=�B���ӗZ�7���/ꗏ[zOD�f���&p��9�a��9tYx\{콜Ȇ��R�/��D��!�h3^�����J������}e^�WT��fH�������\�H��)z��nH1�'��̛c���r����Y+�|-�����j���S۝�.���~��W�%D�$���=三�7����y\� <on(�^&r�+�4�"��=[c�
��/��j%	7"���h k��9�
��^�`X{1L�}�	~bd~���-D���g9�VRÐ�b�^D[5�, ��;}�	ѥ8V��`���{=�������G�\���bhhB^���g���»5��1y�ʦ��hFU�*,���bl��/sE�!����Ih]�����\"�{���YN����)k����ǤuB<U�C����2�C.��W0d<��|f�A������D���O^�"���b:�J�f��f��y���Y��f^�$.T�>��enP�3��ǎ���z�z���G��E�1��fbV]��<?x^y�3r̓ʩ*29˸�7�ځ'@��U���+���dMko)^�Ղ�p��1w@cH��H�{�eĎ�2�Tӫe�B�~<��<`�f|m��h�$NM����h3J�2UI!=��� ���F
���C�̨��<�J{���4q�:F�8B��er�*��g���ͬ�{8|˶|�	3Wc|�+���˼���_�3��ǆ4[��)�D�\��N��9L�����6q\�np�aݫ�I�%�]b���`���m^lO-8�P�k��Y��܎���<L�"T.�cPx&@'Kz����#cc
�u�n��=�±�2ͣX;DK/s�O�&93^�^Zw�v]��vj�T!�=�0�%4K_���y*�τ���f��
^L�_�u����+�p���K�����F��T��cF���|e6bGV2g��k/Ѯ���/W6q�g������I��5�"I��{7�)	4Z}5��#�0�t�H�0ڿ��
Qx�?<���D�EA͈��
����Ӧ��z�JAGc��6�	�,(\���{D�<-,���1`GȺZ�S~�#�J��7|Mb
Q��� ��RI�rS<��P:��.n��`H~+�R�F�%锩�7*��~7�ԩ*r�6�Y���ʼk:�ѣm0[d[v3Ԃ��1{#������[� �c��ZC�MВ���+��9��՗�U<K�Έ=:I�/�g���<�l+h�G������B�CJO�ՌΝ�cI���t ݎ�mc�'������w+r�ǥ�t��1��<f��SS[1��<�I>�|	q�%�KVލ���^�$���CȖ�n�\yI��F��
N�C!�i�B·{�ά���i�+p������B�nw�9d�=��O��_x� ���P�7�yp�P�Z1��q��mW��=���?5h����y����*n/�G�^��h>�D��r��ߏ���\��;��Q/���P�<��-�}��c����0에��x�l�"��+WT��lw9�^+�%�W��?�=qzj��Q��><n�@r[g���#�jكS�';G�0�>>�5��>吷x��8�>�P���#�f��`���C�"���{-�(��o����� /3n��F��Pu@S���M��u���ru��f��E�fFKqsMk8*=��n @8��&PE⧒��G�:�0��7�����Di���Otq��X 8m��/�.'����N\����5Ϯ��J�\yeI �*��8�����U՝d����y��4{m�ԃ�(K�QGCa`�Y�D 3�W�_7��1��a��'W�RNABq� ����aZ���V0�Ʈ���U�oHć��7��M�[=ѓ7�W�P�i����Y�7>�{%2�� *��8.g�v;~��ڧ��dO���g5i���ߑsc��w�\��wuڲο����xH�%�`�/��
���R+�4h�^�Pw����@	��-��{ѭ���k��<�'����t�4*�=���O�k��W���g��qL���u�p�z�А*��H]�!��/���ruJ9e`(�5<��e��u�S,'b�	G�����p�C$�/bQ�ʒ��딏h.�{a!���&�������>���:x��Rǿ���_6��1Oh�݇����|)o?����4���kp��lQ�̘��gWR�$�0A���؁�8�e���ݰ� �ĄcX�6���h����
�.�[���"D239[�꟯{:e�"78��As�y��.t�U�����eN@��3�E�
X���Ǵ�w/�����d|`�լ��\W����_�UV̇h5���ޏX����G!k���}����L-v���|E<����bf��:��bde��g�|ݠ�6(1��<mn��<�uBC`�w#Bf����m�)����ҭ��.�Y~��e���޴�=������m�$�����YF[!� 'r��"<�8�L����k��H�W�e3R��4.ZR��+�cM*Z�g�Iu���+�xV
���;o�-ov�e����J���!��2�Y�;Ή󈯋�/)�E�#�+��	�ul��(Č:W��j�2���Q��Z)Ȃ�Fze>��M�A�)�o�Fi�K�tn�T��C��5��7F=p���m�t�{3�[&���H����/������a�5D�m|h`ޛz|;��t��x�v+�.�u1:sGf	��&wNǥ�[�^�Л��N�Gf^^�v��.كn��o��1���B��{0�&��w�5��qT���gxM�oC�P������]1�'�@)�N郈u����4���@�󌙨�I��w�_`�>���j�L���d}6������H��0�ჵ��M����
�}뾋�N�﬩ ����	��ޕQ��V�FP�P��G�����p���ۘƊ�*�_�<��'N��-��T�̯��!�;�Vׁ�.��B3g����cP����dJ<�M$��x��H�kقb)t}�5�=����s����T@o>E��KPy8��sҧ�%o
b�
¢�?@+��"�7,�P�JY'�]��q��S�B7M��� �+ a�����GD  �px�m�Cq�PU���&�')�����Cst����7dٔ��o�3�~`���<Է��]
.酪=b����S�⅃�y����w9�sF��f׺�h*f�xSD��\��NkmME�� 7+��զ���
�\9_��1�ȣ U��A����f����y�g���+.r�*����3�t౴3V���xl���ț��I���q/R�a%�qM-�^>�B:�]^�/g�A�G-�3�f�<��ٴ�*��ʆ�.��sm&���Q^�6hB{�p,��t�SOοA��Vq�&/K�G�z5s��e�`�+2�M��(�'���]FR��~X�"��E����N���I�e����"ӍKx�>��K��[A�ǩ�n@k��FC�ಳ3
[SHl��jM�L��i%Z�	���h�=!�����|��ٰj�d�|D�����(p󋏻�
�#�M��<��g\򋖎|R�L�Dௌ�y�>��R1���̨O-k]ְ�4�:�\X5��Zhn�1U�k�C7���qOũ�b���0���#�p�����$���^K��6��k��"Sy���_&�]�>���ϔ�1�j��!8�0�%k�n���x,;�$t�@n�~(����� ��y�*�h~�Au�� �Y�]R��60D@�3M�n�M�ϊ�+����?;���J��R(�b�lo��%O��/oa)�L���m�&U5K�ۉHs�8'!�R]]������)n=���dH*Y�(x������ꛢ�m|.^��'ؤ�s)r��,���IEg�v��a�<v'DC'o��4����HW��g�,H�l�~�Y�=��C�B7F��+K��h��>H!vr��7����J�����C퐠B?�«$EK��+c���}���.~���GY�s��]MC��K�}�u�^P�-#��᷻4ɹ{�0P#Vd}��CYb�e��SaLajW��%�hf;� W_�|� |�X��i���@4 ڶ�3�e#Eik�R�K��z��=�y����}����K9�������6�9�mc��N�?�]�qg/8���Y�N�7��������(c���A�w.�JX�6��n@����7	_겪|[@�����Y�%�]GDy^�?�;DE��K=$d5g��Ќ�Y��;�4.�nM�����"��`��vH�4̪�'a������NI[}-)�'�p����^P�4H?纑�v����Ci�2ɋWD��G
�≬�)���Q�_Cu.�'e�%>�9�����V'� �r�1� \v�F�HK�w=)N��P�{O�:�݅ёůs/���8�)g�5I��z����?���%�<�W�]��Uz�،o��(��l��Z�^�B�7eV�H3 g#U�;p��US}��V��w'F��c��.��P�lAx���M�V�J��[����FK[H�<�N�^FH^��R`�X�ھ�>ET��]�����4@��Uu��Uګ�$�u{|�Ho\X9�m���M#��H�������b��5�V�N���'4�I�*^Y
��s�/�Tt״�s�h@"�����>�S�������;~$�y��il��[Ӈ���fZ��U��㩒+l��l�r�\���+�&7(���?y��F�s#��p�=��������C1�� �7rmr�j�����-�}�� C��R�U����d�_w�]��A��� 9���;Vc�YT7[H�R-k����Q��Q�y��,�Z��ﶛ�{D�����*f�jO�_��<<S��+M�8�H�?J@G���k��L�y94��Oh�z�ڍ�ܘ�Q����5����m��m"�}ؚUsu�r]�9��p�u���=b�d�B�t���+��1�c��Т��8E~fb6�A�������P�������� �*4g��T�\��皽D��V�9s�$�5�Ì_q-��: �Nto��L��6o��np�[�^x��<Q�h��"��g5�M��t�k��*�q��_�o1�KiCO�:0Kg�y:{��u���Elu��68���%�=uA�kcT��d��H;�Zs�����e�?��.�<w���hv��+��SEa�N�)��n�C6�U��/HԟK�O;����1	�ot ��GV����j{�-�o�Y����B7�A��NF�[_�F�L˕l�	��C辈
����ꭐ��;�r�_n�9A9�O�U����%Vj�Be�"����y=�p~���bO�	��%,}}F���<ZD�q��2˥��%�jT'����6�8���Uv�m�i���x+ ��ö��z[j��D�dwK��TN�dh��8�s����Q���y��VD�ϕuq���3�iXC��ꀔ�ױ$t�F8�;O�:���?N��
���E,;�/���]��m���Q�o�{3��^�T�5���J�;�a�ܳ��Y����+53�uj�'�7-�Wᆗ"/�Qh�fӆ3�c�1�b��AE7��U��%g]�a�Γ�3E�1ȩ�&�a�hM�&<����]��%�7��~ݿ���RjV3�EEhS������b2�2�ͼ��R� S���Ca��,X�_��L�Nn�.w��
y0������QÎ7ܓd�cm��OF� rF.+BL��H���}��ĝr��F�V:wM,�}̞���){� Ѭ:;���ʍ窕��1�W�GFY�6��2�cӉ�H���,�	��	�#I�C��H���iÙ>��b�۳"R��%��T�Xk�~��oztg`�+uZ��;m��A���}�8��t@c�])2̺��EA&�D� �PB�z��u�&BK^�n����[`�	#2��U�;��8�Z�p�wjQ)%���[9�e��Sv炲l�E�N|D.H��=�~/PX��+��hS3
�C��W�4A����0h�}�s��	I��J�p�vZ�ğ	o��������x92&��a>(�5�gZt�������9�<�8=훲C3��\Eg���
u�8ۂD"�����Xa=1�e|ِ��j��9��N����?6�8%ml�#Z�M�2R��L�h���v�n���$\�����+'	*�I5nK.^���F��r�nU��q����`-<y��Z�o��ԫ�@��.�4�K�^;�K�䤿�-�K!S���PsÞ-�>�>-�q��3֕����&��KG�F�ES<- 6Z
;쓮鸄�:�P�Ŝ�r����M�K�R�';7�x�L������Fy(�;�z���o�TEK= /��^o����h��'ݿ��yB������~�fO�mj��D?����  �\������ЋӇk�3j�d{ ��?���ha�Q�v�*�/��o=��T)#�i"v	$%��$տs��y}bW6�Y�u�:�~	;9 GЧU�H{��0G#�_�_gNE[�:��]ߑc\����,.�(C��zy����9o=�_+�~+��jK�\�V��Uź����!�-Dp]�Fdl8�OKZ��`�ΐ|3�Yy�~j[�Kg�Eb�@őcl�>8P3"�'��׾FX,�]T�x��a�t�,6�倴�EZ�P8n�Js���/���K���4�YJl�A�0�!M� U���u#���պ�Dc#�8�K2a�"�#U���{ꖩ��j"lOä�F�;�xE�=8�z2�Or��B�n���V{��� �S�\e[:���W�	]%��*5�6UQ��@�)
w�XLQ0"P�X/Hᚚ�0ao��J��=�Y_Es��$Y�#M|�wRC��­��2��S�����y�V� ��J^�6���P�Mؙ|3)"�&�zg������\�#�5:|�M`��KE���7���*FCv��%��ü0���8g�00�6Ǒ�ڹ�H�R�7�7\�"��k�����#dr��z�&������&�8eX��q���SʺlB|k\������'� t��
K�_c o���9�k�TTNR�����;�	U#;�~�0�|?r;��y|o�-��~��M����a-+��K�E ��p32�L޲�8� ,ޭd�u���ua���V���>K]�k��e8�Ř�A�<%Z+���b�� �>i��	@���S<.����Z�h��r���*%x�Ey�D��i�I�ѶQ�$����^�lpp�v-UxB�|��i>�(�ꪘ�dS�pY�7S�/}Oͩ�[�%$�C���*�La�fE� |4��H�(�<���KP���,}�4���\�ߕeO�È@��	��4������T �:�ߜOAU̼�',L�ø|Էp9����xq�A��e����k�.��2,�rkQ�;��ȳY?,��r���CUӌƹC_i,���pL�}�/�Ů�bT�V�;�~�mF�j�[+q��T���}�ڷ$����&��fÊ��)��5'��f5H�R5&�X:v�Q$C�z��k�g�TC���*j���wm�S�H�V�e��4�����at���g���,�������1���l��h�d!Q���1s�|9��YP��
������ᄑ�攸���h6
e9��;a��b���IpaՇ���z���ř���]�)����5㌽|܆M����1p��E�aW�R(_:��]�!�ë�)CJ��*�/�����a���^Z�]�N]���F͑f��:�u�����`/?+z��y����C�����y�|���g�2(���E~���*�ݽ\����������Hs��;�8ᶈ���|�D	AeB���O^�t|��g߿�˦d�
��n��� Ѷ��Yu;ME��ug�c[*���P�9@e���Cce#+a��1�zf�p��E��իfs�u~�r�(u��2h��ѧ>��iIA-�0;�fw��V%m��3��=�L��q����
~�����;L�g�!3wD7	���
;�4Xќ*}�Fg�1J5ѿg��]��=T��M��>�GK����������UR�tdJ৉��cb��G�Zz�_^��˄%�1�c�*��%&�l/o�;�%�4V��s��ݷҞ:�\]�/�S��mm/B�}�[S�����GWx���n ��I���@�n��T��ʣ���dbT��[-�'��r8=%�q��ض'oz������!�մ�p������W*KDd�!����|���,�'��4ƫ�Q�̠C��tvwʢ(J}��PƟ�f�c�l�]y��4�����A$��h����8�i\���P��!2�N�
􅷳��u�.[aV?��)m�y3�]������s��45N�����?	K:�L�L��IVj���y \��a�"���'��X�q�c1
�+��k���)L�
�t��ʆc��u_���K?�ϴ��V+�%��
���iL��<P^�<P�r�Y�GPH���-й�S��G����_�k�e/F5��������
����GH�M	̻�����ޚi���_k�R��s���<��K����֒��#�T'&��\y��� � �(�x��Gb�6!~@���0ڱL�QT���ֲ��F�
��.����=�qS�leZ�4�涑��zԠxڂH3�"c����L�&�[Q��G��Q��3�r�"+nH�펝��7�X�!g:~����3����J�����6�y����FX�b���'�o+�;T9��7�l����hU�&c�v���C(��疶�m����s�����jr,�����D�j�Gt��ih^_^`9�w�t�.͆�"k��},�J���d���aw�D�V�H.*L�ԫ�+�1��g8&��l�z	��1/����V�T�tN��P+M)ۈ']E��!�D�̰7J� �̫
m��oI�
�[�eo+�?�[?�*��W�V\�-�}$��h�� �.��9���P��`[�s�� �Ur0I1CB=����)��C=�8�����p�\�Oܷz�f���(�<���E�mm��w�U5���T����C�&��^K���|��J�~ �9�&�ɵv$�G<:��{}{��ɬ�51oL���o�VaE)~m-�p~)�ͬ,�qδq��y�{0m��v�����k-��f�ނ}yY92+�g���E��̥��0���4�x���Q������'*Q�
�Đm.ŗU@��2OpmYۤ��0ܕ��$uX�USѺ8?������B�n��1�w�@l`��ZU}2qQ<���Z�����@;` K�Dh䎵�Lg[�^7�A-�?�on�$\].�������t��u�W�7�rڢGdA��sx:�J�`Rg���2s��� ���ڽ}d�U?*8��#O2������>=~�w�r�e_҉���nR�>���BЮ�X��÷|���`�?r����xx�+�"��RP����*tѢe9��n�T$E=.���V0�O^���oݑ:W�JR��C����S=�ُ�&�7
�YpF�@�F٭ru�º�b� 	G�����"�:���R(�]�����b ŭ���*Ks�6@���H��e�[��|�x�D�r��LLc��DƁ �,���0�mdp��n�*��Epy���?��b$�Wh/�qu~�찲z$o,�����*�QX>T=L9V�;@���o�M���%�IŸ��,f��'��>�QD���H�U�Pi;d��I����.���Fj��׆=�:t�W@�.���-����R�3�q�1"�`]]�����ӊ &��G���\��r��$��>��)-9 :Yџ��.�kZلJ��� �N����^��^�9���ᩏ�[�s��*�z,��ގ�K�5�X��`��w<���'�B�\0���ȍ�|�"pvKc}h���|�,kj�m����R��Ǒ�E~�OB73�x�.B�%�~Y8g|0���H��v�/m@��'k�f]���HF`t�+�xtV�
	e��	mg?��:TN;V۔�/��m���$�>$A����ь��+�ƫP���6�h7K�y��]HΘE���ϽEd�-��$eH}L"h�6������Ryc����ӄ����#�V�Yh�	ph�zZ�PC���%d���X��.��#�����ˊ�և�W�����R�ùQ�>��Y��T�{��@dK��g��}e�(�}�S*#�2ώ[x`�G��o�ڋ����*���K�O�2��V���;� ��+��$����m�7�:�;;�>ג���§�'���5M_Sm���B`x���P5'�|WPTd��.�օ��2���F��ۓ�!{��j���:�n��1<�_�<aD<�D̊���	r�b��E�o��|��ɾ}���J�(�d�:�"��aÅ^oN�O	���nA�~&@B$����t�����m"Y�ǔ��!+S��R�ɒɜ��X:����ϩ��R�[O�4����7�e�p"j���T��}D��$I@����$?(�+\Y��37�>�K#ni�����<z5�|�[<�=���i���-�(����֖�'fX�o����P��w��+;E�Jԍ�&b�J����9$����5��<ɼ>%��*��ӆr��v7=�IThm��9�|ϕDu�j"��@���Ѭ�ΐd��_�Ç-{q�GN�,���@9܏�]/�=��w{��Z��N�R=������N%R����ki�x36O=�{i"kɦ~�=z����N�AQ,ȰKZ�)M�Y�}�_T��
��Y��~9���np�k��1!/�y�����*2������XV�� t6|��+�pZ²�Τ���1��p�C����󴩖"����3/a��=x.a�ZY��&��j1�Χ����:�$J��j�Ȇsi�)	�U��u�~P+� ��Fޫ����`M�� �f��kN �J�8)e�9�{k*Oň��	���� a6?.��9����_C��L�'ӪN=r%�1s�&o\�XZ�a�n�Tuq0LC�����ގ�]9J���`�$�'Ւ�ǻ�殮t&T���\�������kxyQ @����lOs��RZ�����0GXZ䅾0λ٪���i���W�o���+$pk��Y��\K���~g�)ں;��!�����C����Q�N9ɟe���#�J4�o���1>�[K�`�uz��ɴ�P�y9nzxO�EǕ�������z�W�J(��8؊u`���B� �7J�r�4�C�w�nc�>1ūA8w�p?U8��D��b�.�ġQ7�~&��-��>����8F��f��xo�Xڀ�cQ86,#�k�EC<��V���H�u�F��Љ9��%ӥR[/���SyuW�-"{O��tK*���%d"���$���|�ݫ�*+�DaJ�d߼y�U�]t�#ʿU���I��Lqs���	;G�[��u�E����u���n-���	An��ʙ���z-���^.!�ǌ9��Լ ���~�J+�g#/ݍ�U�)�y��� �Q.�O$���G?�\���E��poN��쁑�?��,�Pm�P��$��)����~����,��k�A�r�����7�x����+��d;gtu�<F��9D�[4�M\��i����.�5or�ᴊ�lttM���w�%7rm��%��e��:��%o �ʹ?C��E�T�C8f�A}*�	@��y 1�|H�1��68ϰa��+T��`����%h��gi��*���kSk�sMT�l� �lq�y:�5 V�l9L�E[R��c�ќb�+5Y
�����΢O��q��9M��D
�B
�Y���ĔO�p_�2]�������W�Y֨[,[LՇ��*�P���4�;��ǟ� �P� �٢'��K�/ZH]G��z�3[B|�:Й����=8����M�ϝ*��x5�k����R��8����B�f1�B��Ub����>i�{�07������ZQS`+�����{>x��I��X |[�9YrKFfu�r�u�)�/���!:�:mP-���Ku�0���%%�����d���Q�T6�������Ÿ��]��k�bf����Z��k�)fq��35�Ȱ�)L�ES6�owh��J�7�ݳy�'���U��S��x�l�_a��\F���Ib�T����u�O\(�������G{!�^՟����%��yd��n����h��@��ʑ���ѲM�c]��wD:D�����?uj<+8[�mk*z��_�Xfئ9�)�a��%+�*Y�.CL8�i ΠK��Ͱ��U�q��;hɝ�w��0���\ه,|��E=xcP�AU���*�T	���b�n4�����,�*q/�:
��<�����W�&�A(����?��z��PP{@��'��_�4m�;
5�x@y��X�0��J$����HҾ�*
�k�oן� ˭�9��?�a�,�GM�B(u��!	�R$0ȑ
B�զ�6g��j����o�}CTeEn�S#����˴���v�Cs�s��?�a��E�����@a�Ã���z���B,���#�C�d�̒{�ް ��n.�¡\Q���[ǴL3�����Am���%ǦΦ6`@�b�Z�M�ΈCIB9R��$+Uo�C���������LѴX�KD7�E�I����v�/2�Q�}`�����,ޖ�r�e��N��_���4�%�t����o���Ϡ驹ӎݑ�(�n��$�:�9�4ќ�?�#��;B|��Q�I��m�
ՈHE������h}7_%;���{��il���#�G:�&jY%���L{��<~��(u�I��z�Su����eSSH���Q�g�q���"A$	#�p�ub���NL}?D�k����!b��!��r�97���Ѳ��U�q�T6����<�}�fF�v#�1S2�n�^�A��$8�^h"̂��E���a�����{,�m߶���'�:��3��Nk���Dց����X�E���x�D�:z�MJ�]����J�3"�:���0��;������ѳ.x�BT�2�I��`soJ�����Zr������|R3Yc+�Q��쵯�	�����گw�@���Z����̎���"�OHEʺ�%z�V^��0�)��ns.F��4jHMոZ7>�,�k��/?lF�h�E�`@�NGR+N`,����jn�m�����i<��9�)Ѧ�f����&!�9��_	I����u��A��-�M�j-�2�� �+��X*�9kC�ە�?����y���P�E4�.Y��5����*�������`�
�*2���u�ߐo�ǦQ$���t�WJ�u}��4Ϋ��v%���%[O��$�M�k�cp�<�x�mE#+��$�s�Po��4��jUջ̅9�[��ݤj;�-���r�7���J���XjQqF2��s*�_c����kL�����G	�hF�~���?�����@�l��A33�ȎӾ���ꍽ��K"ߗ
��Q�%r�'��6�Q��bE�l��'y�<���ImeflO�q�O�y���*ܳ�i��l���.D�wmN?�\�R��*Դ�=�UP0����c�$_��bB=ю�*���q�|%휃�j�PWN"�(��^zIj��������Dg9�e�r
�g���B�5\r�<���߈�1���7A`D0ܯJ�4�Gro����1�`Gx����/�����L�n[�B�_t�K���pկ+����b}�FRx-0��L��j�	�Aɹ%�QŔf�w�f�� {Q�Ž�O�%��i��L�}��);i�l���T�  �tWIK�)WD~��x��������dvcf���pXj#�d6�tf�A$rU��ۜ?��(#�=�����ra!C4!������)���)����0��m�