��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�.�&ʺr����$l����<�2�]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPc�k�u�}�|Ѽ�r�ν��e��eG�I�?g�f�SL�<.w[!�� Q鹯e)�Op$=���u��N�w	*D���y&�f��+K��[y��ڂ�Vs>�+��k�:F����/lt�3� P�;��1�-��⫯g*P(�C#<�:z����uP!ߌ��˼�{�&��lV��n��oNaW��4J�Ś��
��H,7f�t�뾌��ߞ�:��L���om�Q*���T�K����Z�e�g�]��s/$W�o?=4��{0��d#m�sj�]:#���c���`�G�YAds£����&����S�BgV�g�0���ή��M�5����J��.���6��H4�
� �AH�}��� �Ȱ��-+�T�8�hF�_!�>>��S�O1����h��]3�;���[=�%�
�R�+�hV�;/=�n;i���2_�q�JX�����@�>��+R���RL�a)=�y�~ ���������ߤ����Q�=�>�v�ֹY���8＀�L��q�Jp� ��g������a6���r<����}�a
��{0��d#��翑��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A����2�P`��������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW�{b�2"���Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ�^��+o��sKJ�lق�����'SR����.�}|��ι%9T��7���S5H�j.F�YZY0@ìOd��q�G�+��T��`	��
�+����/�!��-`���[ b�����,\ަ�It�-;O��M�����$��q����-���լR���*F�57�@��+�wD~�	��4s�ٷ��M��o���hW���1�>�&����1~�u�pჳ�e����te.T��A��N���C�vC/�ɨ�-�}���ԯ��X��a��X�Ϲ�x���{i�etxUU�Y��N�0�/<~�a_0y�'W'}�����3����LoL;wi6�Z#���t�|̸9�7=���������qθ
��xY{^@?8X�,x7�T�٥��T ���'��;R!�#��z�mgI�9����'*`�lChg���z���Ȥ,��/����U���hNJ�p_��I�����7:�F���2�EN�@���k�� ���3�ҺIÙ=�Hr��~-���I�R���F��c��Z��}��	�d�bzP#�-������4Q��#��w21�X��|�C#/<���q��!�u�ǭ��k��?��}��7Q�� +@����������'�=�OT���0�4z�S4ٗG�D:�]��H/!�S�av>�)'l:}��Q�Ȩ�+)	Y���
Ta�~�4�k�|L����ҭٕ!! �ָ3�o�:��o�Y�#�Ez��R�>}1�l+Tf]�i�#�l�-Px���H��U��p騥%�W,��{���7K��;������(�\���W/�������m��Z�
b�tU��֜��3��TG���PIÙ=�H�c��Э|;>bv�E��5�F��������5	���]���c�A�L'�������W��_�ړ8���/��4��}�<�N컽kg����|g�Y�'���Xw�j�7����'�e���"j���b7|#9���Y��
�iC�E����F��j��\w��0]%��C���+�
�c�~��j��\w��0]��0�&�ͭ�E����F��j��\w��0]{k�h�+m��q'��7G#+�Ǘ0z�cUL
 '&1���D���J��8���/���:��ӰӒ1�:�Ω�P�p^��J���t��.�z,y�%���E�EYZ/�矘��-n��I�?g�fWg�X1����5y�$����<�2�K��3i~���u��wb�S��V��(8�q��Z�y��s��3޴+����cG 7���9Ի0��V�0�!�&�*�p6�!"`�P���$����Zh"?����ǁ�D=��]ݸ�.�8K���iM0�3gf�z�;qǙ�d��hw���gۮBez����AmY�f�4 T���&�]�F����M��_(����@҄���G�۰��{�w����>s.���b9���.M�"��Ӗw�c*����Xa�R�+�_����=k�Rm��̬��[�]��z���;�A�Y	���^�^�� ��͌U8r��<���E�=��ل�9QHll�nf�O�ˎ�����`�N�hX�0�/�zU�=�����?*��.��6�^�� ��͌����҅�#��3���Ct�w#��@#��`*���0u�\k|��.iA�?^�Fa���d��ݫ�Q�n=j��E(%����������iM0�3��w�nV�f�	��8�##;�:E��$vi�N;=��c8?-+eN��zʛʑS��_���!+}$|~ïSup�xg�����{���ض�Ů���zPt� ���1#��Z�����XP���G�@[E�Bn�*5H8P�@<>��%�}L�@��J'�!�5�Zv]�kk�cP��л�+U�HJ�h4�9B�K��\�v�{=J�����?���^�����=j������{�Z���!s9�L���hKR�wX�� N��r*�1W�V�bS�-�=q�:Gz�LQ �� 
~�F���r?j��69Q4���x��W B��A=�� �C� ��Hځix�&Ofۢ��%P���X��T۳�͕��4uB�����ڔ�f�uojr쇤m�O��Ü�/�zU�=�����?��Si�9�׏�����M�~���i�x˗9��6�8�d^�ϓ�Ü�E���J��K�MJJ�Y6�B�n=j��E(;�ѽi�|�0��GP���%��]��}R���rѕ���!�_$!�e����ɬc��WN��&��w�+Y��b9@�g��l�7L���o�0�[X�b\gXA�d�7�W�l��9�vL"\�$Ǜ�?�d4)�\��L�D2����W�럸���c�7*E��|e��]�!�����=�߼
�dA#�V�Y����	�_ȡzab����j7��i�j��~�3�Z�I��(^,��]p+_[�.���e��^��q6\�����4�M����`,�"Ũ����X�"LT߫�%�$�
_���Ȇ��S*��Ֆi�8�O��=�"�Z�p�����[�������C Ln��S�W�.�p�2�zgf�z�;qǙ�d��hw�K-��V�Z$�mo�6L�J'�!�5�����T��z~��x?���Լ����R��c8?-+eNy+�>K�VE�g�;�b� �4�r6�h}�L00:�b9����'0Ѵ��V����aU�`�K-��Cҷ��e,���D�MJJ�Y6�B�����6���'�e���ъ����K(�
�cc�V�{���G��R���c&;O7}�»1#��Z�����XP���G�@[E�Bn�*5H8P�u��0��4��
�cc�V�AmY�f�^W��.P5 ���V�Z-�B��cȬߝ��v�2(t��4l��z��_#Ԡ/����KQ�D���Q��Y����LDπ���w�nV�f�	��8�#@��5P���\�}^A�T�g�v�!�����uG`�_BI�-���6%���UbG��V�6IWJE�r���秹�3I^�vKw����qc�U_�+X���=ў@'���Xw�j�7���c8?-+eN�CyW�f�tR�wX�Ռ�O;���9J\�e
`�}R�򳄖�|����=%+]Bo�A;h�F�sZ��;ӹ*"v%)��Qcm h�]�!��	Ǹ�y85�-�)�{�Z��s��R�wX����?�m�����x���y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL�ݵj�<oU��֜��3�T�\ ��W���g
�4�C�w:h���_��*`Dg�8�Hk��|��-Wl���[w�4��<Ր���hn�����aUyR�b!������16X���p+��]��CJ�dR�wX����K�Q�+�4�i iJa��������ܖAA/���G�c~C�|��m=�L|Dt �PW��a��K�TR"K�g��U-�e(��w��x�ȳ�5�(�T�\ ���|.�Tӏ7U We��M�1��n��FR���'S/�_wπ>���9J\�e
`�q���ʭ�O7}�»����Ck�MN�3�Q�D��̣����F�z�C���#�^�&F��C�s��e�������hM��1o�l�P:�R����s�N���IQנF���ϸ�U��?���D|	�õ��Mn�;��c���XyR�b!����`y���pzl��a�8���SY�N iJa��������ܖA���ol��t�c~C�|��m=�L|Dt����U�#y �Ac�N�A���1#%�"MN�3��cSS�b�(Q6D����z�C���qg2�K?\?��~]l�*`Dg�8�Hk��|���DD[w�4��<բ�]Z�Cď��/V�h}�L00:�g��U-�e(��w��x��-��U���T�\ ���|.�TӏpR���Ny	|4�F�(�X)󿥠&���Z02{�"��}�u4��d�bR�wX����K�Q��Jq�Y���̓q�i&.`�]`�?���� ����C �Q��Y����Qs����[�=�5x�9B��2�_�d`:�qP�㎏qló��U��?��]�W�m��8���/�a'�<� \��2{U	fPߑ���K��Q]� _�rs�i�ק)"�僁�cSS�b�YG���R�wX����K�QڱA�e!�.͌FE�K�7s�9���o��S8��A��H�cBh}�L00:C?�Q䨈�z�C���\�#$�ÙAx�:$�ջ�ﻋ-���>��l%i�-�s��d�\�F萡x��t/�(�P╳x�X�"��l��{N|3�cSS�b�i'��s�e|q��M���Lu�>�� ��6h���v�䩲$���5�R�̺l��vC�|1,'����0�zG��"Όd)���M7<Q�D,#�`j�cSS�b�YG����dh_��tCdN�<@Iv��nt=:�b?0s��0�ʂ�j�Ï��	�l�lM�3 �[�{3^��=�O�-v�*_�mS8<�n8"25V��O@ Tߌ�\�����aU˙����Wѫ���Uh1�P����v�\�w�0i%{�"��}ϻ�_��4���܂�����TS4�04�jf���F��O�<�P�����os�鮊�����n�Z6j�"Hs][.6h3(_6���Yx-�'�b�  �ҋ�;Y���D���!�'��أͽgF"?���p+���"M�RZ�y��K�ݽ��������D5�|أͽgF"?���p+���"M�RZ�xkx U�_@���U���&0�]̽Cl�;��|B���8U����_��*`Dg�8�Hk��|��m�d�6���!�=�ߝ��v�6t#f���	��"X��[�-�Vb� �[�̷��3h�/���k��Q�D�䀄8h�Y�Ȫꤊ�u�܎����~�֢);�A�T�g�v��o
���^��"�C�˂j}�C���&��vt������=:9��Y/7 �4�r6��cU�tF�"�S��rN��t"O]=��Y�$��b�H�������p+��i�~͜b
BqBé��U��֜��3���HK�A��n� _J�/Td@��c�����M�~��~@�H@'X35Y��Ap��E&���?�d���&���Gh�d��''�|7�=N;]%z���5��Z"��a�d�yH	Z���/:���lC��U�T�\ ��.��惏�''�|7�=N;]%z���5��Z"ц�U�p��1��C���5�%]���a(􆿳�e�&���6�a��T� iJa��������ܖAA/���Gx�p��F�A�T�g�v�"j���b7T�K�^d��ȹ� �tw iJa��������ܖA���ol��t���������*����6��	���`y���Ż�&ǥ��?�d���&�!�2����|��G�Ȧj�Q�ͼ���ݼ�:zWN�c���Ņ]g����ݰ��W�.R�ix`��T�$^(?��"�SΣ�S�x<�K�'ž1�|�'����nyֽ'����}v�e�q_҂T�q��n"��
l�Q�D���AƖX�y���?~f|��d����̄$Sgbd)H;��c���X���%���@f	2J������_��*`Dg�8�Hk��|��!�x������p�1e��0�U+�qbp@�*���?�HKM�1��n��FR���'S/�_wπ>��M��b_X�XV�b�z'hۉ)��R��삍(�V�ܼ�l+��H����ݾ-/�P��f��T/��k
+u����g�Z��3��a���!@�f")%n§z'�zy�}�6f&rG��Hbr��������J�j��+C�>��r?j����K�TR"K{H�3)-��Ǌjj�����o�����mbh�O7}�»ԯ�J'>c�~�1�|2�''�|7�=N;]%z���5��Z"!�%2��N�� ���E�����_��*`Dg�8�Hk��|��m�d�6���:Vg������ �}-�п� W��$0���>�����nR�N�o�y�<�J��`�{CE���'!msR�����נp�Qe�L�D٪������&^����_�'G
��T���xvW'��}�B�����׏�����M/X*F���&�2Ƣ�IX0F�M�~s\�̻W<u�g-�U��)��h�ߨ��4+©��.DR�&��b����&e*!�Hѷ���A��$�Qu���Lw]�D���z?7`8ȵ�ixUS�����*��|>����n�������+U�HJ�h�,3�Hs8�}�����:P"G�wk�
c�J>w�#Z��s��R�wX�Շ��������-f/]������sT�@�3𗸟�am� W�����o�Ъ���ll�K#4�rq�B�3�B�����������>7�Y�r���	 f�b�H��<�C_�,���� �Ac�N�A乏�-���/�ciJ�B��A=��D1��4���Ut�\��`��t����@|�)��8���e���a-6�DaHP%���e�Hĝ$�pi�9a�Fc��]���#�0����x ѻ��3qV�	PcM�9S����q��k��\�v�07�����_M�<TC���qyJT��rW��]��C ����X8��8���/���K�����aٔ^?���w:&��}w"�5 �Ac�N�AO%^�p�c�g��U-�e�´��'�)�Բc*�r#�ӑ�{��|M1�9$[{^��o|����"X��[l-���}���q%�����Mg.6�kT۳�͕��i1n�6P��4,�Q����W��'�)�Բcf�x�HZ�, ���q3HL�1p/-��}-���NHRxF� l�f~,q��M'�b�	�)�.�ij0���!{�"��}n�m!t%qa(􆿳��ύ�>� ']v1�_ُ�&��b���/Q����ߝ��v�Y/�ܜ�������#oM.�����a�x���Jq�Y���y-T�OB �4�r6�h}�L00:� ^M'��k/��m#'�a[μ3z� �z�Ep�-a�D͢q��`�L]Ć[�_ijsrCm�kp�z����'���Xw�j�7�� �X��E=r4�ё�{ѧͿS����w,��I��KO8���	�)�.�i�WB|Oݤ{!�
ܯ�Z��"L?��پ9�d�L�ڱA�e!�.Y�+�����"Όd)��d���T��jsrCm�k(%�ar�s8��b�Bϱ���2�b=�������AԢ�a\�	PcM�9S����q��k��\�v�07�����_M�<TC�}�����:(���27:����aٔ^?���w:&��ˮ�t�s�'�)�Բc*�r#�ӑ���?O�y	�?�\�
-�:��KY�[b%Ɨ����н�!]0{ɽ�����$��ރ'�)�Բcf�x�HZ�S]�*
�]v1�_ُò������?O�y	�)�x�.#P�j2E�? �X��E=r5J�Ӝ$����b�Bϱ�B����iZ����q��k�P"G�wk��v0�%��U�����zyN'�a[μ3z� �z�Ep�-a�D͢q��`�L��F\�l&�c%=�)�]�!��	Ǹ�y85��C�%����ۯ�����Z��/��\�w�0i%(ξv�釰 �X��E=r�����Z*V�M��nD#k�˟ܒ�o|k�LbfF�5.]��۪	�}a�IX0F�Mұ�*ȣ����W�`�f�cKݸ){�"��}����@����p+����g�I��e�2�=Y��>{�i�C��-�RfJ�J|[��alD�� {Z���ڨ|����.�e��U4��\��P�%�+ Ixcw���Z�����S��C����B)|D/[f^���;��c���X K�D��t䃦�=���>��ڷ�y؛�"�'����"O��1h>E}#���Z��E{'��p���qU��r|]��� a⣃_BO������k:͋��C8�oFJ�u�S�c�7�i�2�L���)�J�I�)�z�����]���I����+��C#�K�"a��ُ�S���v�?�����s�cki`:Gu{�F�ï�y'Ƶ�s0��J�dG3;�hs���p+�����FL�V�8���/�&k@C�Ɨ0z�cUL��G'T�$6$�s�N�|���]k�H��'!msR������lʛ�����}w"�5O7}�»�E�0#�4j�T�\ ��ه� �4�<��Jq�Y���y-T�OB �4�r6��cU�tFZQDu����-�Vb� �Z鎬�������(�����I C�s��e�������hM��1o�l�P��+�����������m�۶t���������#oM��:<��j�P�++�hW�w��fD֌�J8`ϣ6�}"y��7.�O^�kO`,Q�D������B#�v��~ a⣃_BO������k:͋��C8�oFJ�u�S�c�7�i�2�L���)�J�I�)�z�����]���I����+��C#�K�"a��ُ�S���v�?�����s�cki`:Gu{qĝ�&������w:&��}w"�5O7}�»p�[k����Cҷ��e̷_��yC��S8�k��m�ݧ�H7
�߀�}-�п� W��$0���>���ˍ���AD��/���k��Q�D������X8��8���/�n�Ҡ8P  a�o$���w�)>B:�Z�m�۶t�����D�P�E6�n)Pf�� '���Xw�j�7��֏j��[�*5���@*`Dg�8�Hk��|��!�x�����!�=�ߝ��vԩ �E�p��"X��[˹�H٫!��G�Ȧj�E��g�Hb��B���%2�����Vcڗ�q�j�I�=H%�_[X"�T��>C⣔���t��W��-��U����,KI�$�}��w�}�2v"]U����`h��}� �`NZ��Vܟ=�a~\C�~��/�4�ooG��e!�nwUSc�!{p85��:�"�D��qU��rbA���݋Fs��u�x�9��_r/��(��ڍ�-��U��?�d���&�]�0^ݵT"�1?'����!���5�Nn�25����#h}�L00:u���Y`i�7�Ϛ�.'Ƶ�s0��J�d�,e"75�EZ��s��rN��t"O]��!���c�A�L'@fU�X?0I"�`�it�M��f����_��*`Dg�8�Hk��|�I����Q�D��8߄���*t �4�r6��cU�tF���p+����;�),�8���/����-CC���z��n�Ҡ8P  a�o$���w�E���s��U��֜��3�T�\ �͊�51�X�c�rs�i��]S���D[�l��a[�S�� ��|`/+ iJa��������ܖA���ol��t����aUF�7'HR9q�}w"�5O7}�»l�2vh�1�{�Y��a(􆿳��˜T�Ԕ�m��'A>g4�����ρ�@b���ѰQ{�Nj�t<78]�D� nqҺ�Ib��SfȂS�Z�����D�p�"$J��l�H��9�����L8h��l�"!��<63tI�w�g�ˇ�Q��F^�c�����M�~�Y�5� a��2�����Vc�{b�'���Lx�ƺ�M���	�n��XU���#fhr��y�ڔ�.������������/�LBgh�c,q������z�.���f%%eo���sp%�j����P"G�wk��%R[�]db6ڏ� �7.�O��S}o�"_�cSS�b垊*��䮻E�&�y+B����iZ�1T棗���m��'A>�g��U-�e"�A��"�Y�{'%s��v�9˞�g��+˘\59:��lJ�ſ@,�$�}-�п� W��$0���>���˰��0������:UkG3;�hs���p+��v W���}q�!D�t
���"X��[��h�C��hA�T�g�v�i��Z�qĝ�&���w9Z� 0�����*��|>����n�T�K�^d��]�!��	Ǹ�y85���]��^������.'�L����^�7�Y\�� =N;]%z���5��Z"�'��G�<���,Y#A	u�e�2�?�m�۶�so����O7}�»�QNȮ���k/��m#�J'�!���=�@q��u���"6ޭ<:�&.am� W�����H��6�Br���N%'tF��;���R��C� �Y��#_1�|.�~� �����$�\՛��2�k�S�{ �d�*��M�,4#�rQ����(��t�;��|B^nl3Υ$���G�Ȧj�Q�ͼ�����l_��F�h�76AyW��㜿�k���<^&!!HYx����Rd݉'~�zM����!Mr�J�M�
9E��O d�?�ykk)��T�<�Fs��u8�RX7���#g�k��9����4`-7i�J١��ߝ��v�Y/�ܜ���}��9��z���FY�g��U-�e�c8?-+eN;�\��	�8���SY�N iJa��������ܖAA/���G����aU�D�mD�VOR�)���$~�ߝ��v�Y/�ܜ�������#oM������c�����M�~��4e62A�I����Oݷ �*$�8�RX7���#g�k��9����4`-7i�J١��ߝ��v�Y/�ܜ���}��9��z���FY�g��U-�e�c8?-+eN;�\��	�8���SY�N iJa��������ܖA���ol��t����aU�D�mD�VOR�)���$~�ߝ��v�Y/�ܜ�������#oM������c�����M�~��"�l�7%����,�ǰ�͕e���M�@�,�#�j��$P����w)���r?j��h}�L00:;��|Bx R��u��X�趈�w�⽒�;��c���X8�RX7���#g�k��BgG\���De�<[X���H�V�!\��:��1�R��j}�C���&��vt������=:9��Y/7 �4�r6�h}�L00:)�/����Cҷ��e9f2Pih{q��t�3��/���k���cSS�b�l2�_�V��T�\ �ͭNjX�U�6j�"Hs`\��45��wٺ�}aG�k.9Z����t�h��E�&�y+�1�R��j}�C���&��vt������m`%e�I��m��'A>��"X��[�-�Vb� ��1�R��j}�C���&��vt�*��]�3ྯ�;ܙ�c8?-+eN�CyW�f�tR�wX���P�++�hW�w��fD"#��^�D1����,�ǰ�Bί}\Q;��8qV��	��yf��j]/�f� ��T�S���Ev�#+���ÃI���c�90��q�	_����+�^�N���5��x�>�+X�M?��y�if�ً%�^��c���|��RCc��P�f�e�B��6�I�h�S-^^B;�֙�K�J��G{����c�cSS�b���iqj�3��ʄ��!?��~]l�*`Dg�8�Hk��|��!�x������p�1e��0�U+�qbp@�p�-a�D͢��&�j��y����\�&^�����:9g�N�/��dc�@c�����hW�t!:�
����' �^ ���LQ�/8n
V~$�.����hq_҂T�q��n"��
l��cSS�b�ԯ�J'>cI��@%B��qĖ7v�q�8�T�����P��:'���e2o���wu6���ξ�|��U>�f&��'!msR������K�=p�-�	� �~�9rF�؀ǏU�e��FR���'S/�_wπ>jzT�;D����kƢ*NfF�5.]��r�9�7��p�-a�D͢��&�j�ѹ6:�j��5ߧE4����u����Q5��5��φ��<�6�*'頭�Vӗ�e����6�ޤ[QG�